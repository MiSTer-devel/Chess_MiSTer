library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_white_rook_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_white_rook_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"2A000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"35000000",
      x"13000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"2A000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"2A000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"35000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"34000000",
      x"2A000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"45000000",
      x"D1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"E2000000",
      x"C0000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"45000000",
      x"D1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"D1000000",
      x"45000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"C0000000",
      x"E2000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"E1000000",
      x"D1000000",
      x"45000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"65000000",
      x"F4000000",
      x"FF060606",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF191919",
      x"FF050505",
      x"FF000000",
      x"00000000",
      x"02000000",
      x"02000000",
      x"04000000",
      x"66000000",
      x"F4000000",
      x"FF060606",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF060606",
      x"F4000000",
      x"66000000",
      x"04000000",
      x"02000000",
      x"02000000",
      x"00000000",
      x"FF000000",
      x"FF050505",
      x"FF191919",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF060606",
      x"F4000000",
      x"65000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"65000000",
      x"F4000000",
      x"FF2E2E2E",
      x"FFC9C9C9",
      x"FFCACACA",
      x"FFB4B4B4",
      x"FF292929",
      x"FF000000",
      x"5F000000",
      x"65000000",
      x"65000000",
      x"66000000",
      x"A4000000",
      x"F9000000",
      x"FF2E2E2E",
      x"FFC9C9C9",
      x"FFCACACA",
      x"FFCACACA",
      x"FFC9C9C9",
      x"FF2D2D2D",
      x"F9000000",
      x"A4000000",
      x"66000000",
      x"65000000",
      x"65000000",
      x"5F000000",
      x"FF000000",
      x"FF292929",
      x"FFB4B4B4",
      x"FFCACACA",
      x"FFC9C9C9",
      x"FF2D2D2D",
      x"F4000000",
      x"65000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"65000000",
      x"F4000000",
      x"FF393939",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFE2E2E2",
      x"FF373737",
      x"FE000000",
      x"F4000000",
      x"F4000000",
      x"F4000000",
      x"F4000000",
      x"F9000000",
      x"FE000000",
      x"FF383838",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF383838",
      x"FE000000",
      x"F9000000",
      x"F4000000",
      x"F4000000",
      x"F4000000",
      x"F4000000",
      x"FE000000",
      x"FF373737",
      x"FFE2E2E2",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FF393939",
      x"F4000000",
      x"65000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"65000000",
      x"F4000000",
      x"FF393939",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFF5F5F5",
      x"FF858585",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF383838",
      x"FFA7A7A7",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFA7A7A7",
      x"FF383838",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF848484",
      x"FFF5F5F5",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FF393939",
      x"F4000000",
      x"65000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"65000000",
      x"F4000000",
      x"FF393939",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FF393939",
      x"F4000000",
      x"65000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"65000000",
      x"F4000000",
      x"FF3A3A3A",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF3A3A3A",
      x"F4000000",
      x"65000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"64000000",
      x"F4000000",
      x"FF000000",
      x"FF030303",
      x"FF0A0A0A",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0A0A0A",
      x"FF030303",
      x"FF000000",
      x"F3000000",
      x"63000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2B000000",
      x"BF000000",
      x"FE000000",
      x"FF101010",
      x"FF767676",
      x"FF9C9C9C",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9A9A9A",
      x"FF9C9C9C",
      x"FF757575",
      x"FF101010",
      x"FF000000",
      x"BE000000",
      x"28000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"1A000000",
      x"C1000000",
      x"FE020202",
      x"FF282828",
      x"FFE7E7E7",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFE7E7E7",
      x"FF282828",
      x"FF030303",
      x"C1000000",
      x"1A000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"19000000",
      x"C0000000",
      x"FD000000",
      x"FF282828",
      x"FFBABABA",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFC6C6C6",
      x"FFBABABA",
      x"FF282828",
      x"FD000000",
      x"C0000000",
      x"19000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"31000000",
      x"C7000000",
      x"FF020202",
      x"FF2B2B2B",
      x"FF616161",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF646464",
      x"FF616161",
      x"FF2B2B2B",
      x"FF020202",
      x"C7000000",
      x"31000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"72000000",
      x"FF020202",
      x"FF626262",
      x"FFEAEAEA",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFEAEAEA",
      x"FF626262",
      x"FF020202",
      x"72000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF646464",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF646464",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"66000000",
      x"FF000000",
      x"FF141414",
      x"FF333333",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF363636",
      x"FF333333",
      x"FF151515",
      x"FF000000",
      x"66000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"AD000000",
      x"FF030303",
      x"FF474747",
      x"FF929292",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF929292",
      x"FF474747",
      x"FF030303",
      x"AD000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"50000000",
      x"EB000000",
      x"FF191919",
      x"FFBCBCBC",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFBCBCBC",
      x"FF191919",
      x"EB000000",
      x"50000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2C000000",
      x"C4000000",
      x"FE000000",
      x"FF282828",
      x"FF929292",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF959595",
      x"FF929292",
      x"FF282828",
      x"FE000000",
      x"C4000000",
      x"2C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"F0000000",
      x"FF000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"FE000000",
      x"F0000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF121212",
      x"FF4E4E4E",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF585858",
      x"FF4E4E4E",
      x"FF121212",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF333333",
      x"FFD6D6D6",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFF2F2F2",
      x"FFD6D6D6",
      x"FF333333",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF363636",
      x"FFE2E2E2",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE2E2E2",
      x"FF363636",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1E000000",
      x"35000000",
      x"34000000",
      x"31000000",
      x"FF000000",
      x"FF292929",
      x"FFB4B4B4",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFCACACA",
      x"FFB4B4B4",
      x"FF292929",
      x"FF000000",
      x"31000000",
      x"34000000",
      x"35000000",
      x"1E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1E000000",
      x"B7000000",
      x"E1000000",
      x"E1000000",
      x"DF000000",
      x"FF000000",
      x"FF050505",
      x"FF191919",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF191919",
      x"FF050505",
      x"FF000000",
      x"DF000000",
      x"E1000000",
      x"E1000000",
      x"B7000000",
      x"1D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"36000000",
      x"E1000000",
      x"FF030303",
      x"FF171717",
      x"FF1D1D1D",
      x"FF1C1C1C",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF181818",
      x"FF1C1C1C",
      x"FF1D1D1D",
      x"FF171717",
      x"FF030303",
      x"E1000000",
      x"36000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"35000000",
      x"E1000000",
      x"FF171717",
      x"FFA1A1A1",
      x"FFCACACA",
      x"FFC8C8C8",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC0C0C0",
      x"FFC8C8C8",
      x"FFCACACA",
      x"FFA1A1A1",
      x"FF171717",
      x"E1000000",
      x"35000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"35000000",
      x"E1000000",
      x"FF1F1F1F",
      x"FFCDCDCD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCDCDCD",
      x"FF1F1F1F",
      x"E1000000",
      x"35000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"34000000",
      x"E1000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"E1000000",
      x"34000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"19000000",
      x"A2000000",
      x"CB000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CB000000",
      x"A3000000",
      x"19000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"12000000",
      x"1E000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1E000000",
      x"12000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
