library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_black_queen_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_black_queen_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"1A000000",
      x"34000000",
      x"34000000",
      x"1A000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"2F000000",
      x"1C000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"44000000",
      x"C0000000",
      x"F3000000",
      x"F3000000",
      x"BF000000",
      x"43000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"49000000",
      x"C4000000",
      x"DD000000",
      x"D6000000",
      x"74000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"E7000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"E6000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"34000000",
      x"5C000000",
      x"1F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"25000000",
      x"D3000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"FF000000",
      x"74000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"4F000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"4E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"14000000",
      x"A6000000",
      x"FF000000",
      x"FF000000",
      x"F4000000",
      x"76000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"67000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"D6000000",
      x"1C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"4A000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"49000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"A0000000",
      x"FE000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"E9000000",
      x"39000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"8C000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"DD000000",
      x"2F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"E5000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"E5000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"29000000",
      x"DB000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"80000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"19000000",
      x"33000000",
      x"34000000",
      x"1B000000",
      x"04000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"4F000000",
      x"FA000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C3000000",
      x"12000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"36000000",
      x"D8000000",
      x"FB000000",
      x"FB000000",
      x"D8000000",
      x"36000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"29000000",
      x"DB000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"80000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"04000000",
      x"1B000000",
      x"34000000",
      x"33000000",
      x"19000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"50000000",
      x"C2000000",
      x"F1000000",
      x"F3000000",
      x"C0000000",
      x"4C000000",
      x"04000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"15000000",
      x"A7000000",
      x"F9000000",
      x"FF000000",
      x"FF000000",
      x"D3000000",
      x"49000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"3F000000",
      x"E1000000",
      x"E1000000",
      x"3F000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"9F000000",
      x"FE000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"E9000000",
      x"39000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"04000000",
      x"4C000000",
      x"C0000000",
      x"F3000000",
      x"F1000000",
      x"C2000000",
      x"4F000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2E000000",
      x"D5000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"C0000000",
      x"1B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"15000000",
      x"4A000000",
      x"FE000000",
      x"B4000000",
      x"2A000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3B000000",
      x"E4000000",
      x"E4000000",
      x"3B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"14000000",
      x"A5000000",
      x"FF000000",
      x"FE000000",
      x"F4000000",
      x"75000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1B000000",
      x"C0000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"D5000000",
      x"2D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"59000000",
      x"F2000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F2000000",
      x"33000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"C6000000",
      x"1B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"58000000",
      x"F1000000",
      x"F1000000",
      x"58000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"A8000000",
      x"FE000000",
      x"1A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"33000000",
      x"F2000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F2000000",
      x"59000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"58000000",
      x"F1000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F1000000",
      x"33000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"F6000000",
      x"4A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"76000000",
      x"F7000000",
      x"F7000000",
      x"76000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"28000000",
      x"DE000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"33000000",
      x"F1000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F1000000",
      x"58000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2A000000",
      x"DE000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C1000000",
      x"18000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"B7000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0A000000",
      x"97000000",
      x"FD000000",
      x"FD000000",
      x"97000000",
      x"0A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"72000000",
      x"FE000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"19000000",
      x"C2000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"DD000000",
      x"29000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"54000000",
      x"DE000000",
      x"F1000000",
      x"F6000000",
      x"F4000000",
      x"67000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FE000000",
      x"FF000000",
      x"29000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"12000000",
      x"B3000000",
      x"FF000000",
      x"FF000000",
      x"B3000000",
      x"12000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"E8000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"67000000",
      x"F4000000",
      x"F6000000",
      x"F1000000",
      x"DD000000",
      x"54000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2A000000",
      x"56000000",
      x"78000000",
      x"FA000000",
      x"95000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"A0000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"21000000",
      x"D1000000",
      x"FF000000",
      x"FF000000",
      x"D1000000",
      x"21000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"6D000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"95000000",
      x"FA000000",
      x"78000000",
      x"56000000",
      x"29000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"07000000",
      x"FF000000",
      x"F2000000",
      x"3E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"DA000000",
      x"2B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"32000000",
      x"F0000000",
      x"FF000000",
      x"FF000000",
      x"F1000000",
      x"32000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"14000000",
      x"C8000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3E000000",
      x"F2000000",
      x"FF000000",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"DC000000",
      x"FF000000",
      x"D8000000",
      x"10000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F4000000",
      x"63000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"4E000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"4E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"4E000000",
      x"EC000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"10000000",
      x"D8000000",
      x"FF000000",
      x"DC000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"A4000000",
      x"FF000000",
      x"FF000000",
      x"97000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FD000000",
      x"A2000000",
      x"0E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"90000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"90000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"8C000000",
      x"FA000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"97000000",
      x"FF000000",
      x"FF000000",
      x"A4000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"6B000000",
      x"FF000000",
      x"FE000000",
      x"EC000000",
      x"4F000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"DD000000",
      x"27000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"D5000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"D5000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1E000000",
      x"C9000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"50000000",
      x"EC000000",
      x"FE000000",
      x"FF000000",
      x"6B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3D000000",
      x"FD000000",
      x"FF000000",
      x"FE000000",
      x"B4000000",
      x"15000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"64000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"4C000000",
      x"FD000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"15000000",
      x"B4000000",
      x"FE000000",
      x"FF000000",
      x"FD000000",
      x"3D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2E000000",
      x"EA000000",
      x"FF000000",
      x"FE000000",
      x"F5000000",
      x"70000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"DB000000",
      x"07000000",
      x"00000000",
      x"49000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"49000000",
      x"00000000",
      x"00000000",
      x"C0000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"6F000000",
      x"F5000000",
      x"FF000000",
      x"FF000000",
      x"EA000000",
      x"2F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"21000000",
      x"D0000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"F1000000",
      x"30000000",
      x"00000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"5C000000",
      x"00000000",
      x"8E000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"8E000000",
      x"00000000",
      x"40000000",
      x"FD000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"00000000",
      x"30000000",
      x"F1000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"D0000000",
      x"21000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"B7000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C6000000",
      x"0F000000",
      x"00000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C3000000",
      x"09000000",
      x"C3000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C3000000",
      x"07000000",
      x"B6000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"00000000",
      x"0F000000",
      x"C6000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"B7000000",
      x"13000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"A0000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F3000000",
      x"6D000000",
      x"05000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"E5000000",
      x"56000000",
      x"D3000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"D2000000",
      x"4E000000",
      x"E1000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"05000000",
      x"6D000000",
      x"F3000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"A0000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"07000000",
      x"85000000",
      x"FA000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"CF000000",
      x"1B000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F6000000",
      x"B2000000",
      x"E9000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"E9000000",
      x"AB000000",
      x"F5000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"1B000000",
      x"CE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FA000000",
      x"85000000",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"6A000000",
      x"F5000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"82000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"FB000000",
      x"FD000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FD000000",
      x"F9000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"82000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F5000000",
      x"6A000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"51000000",
      x"EF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"F8000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"F8000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"EF000000",
      x"51000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3A000000",
      x"E3000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"E3000000",
      x"3A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"21000000",
      x"D5000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"D5000000",
      x"20000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0A000000",
      x"CA000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"CA000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"B7000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"B5000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"55000000",
      x"F7000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"F7000000",
      x"54000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"85000000",
      x"F0000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"EF000000",
      x"84000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0E000000",
      x"89000000",
      x"F8000000",
      x"FF000000",
      x"FF000000",
      x"FF111111",
      x"FF353535",
      x"FF565656",
      x"FF717171",
      x"FF888888",
      x"FF979797",
      x"FFA7A7A7",
      x"FFB5B5B5",
      x"FFC1C1C1",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC1C1C1",
      x"FFB5B5B5",
      x"FFA7A7A7",
      x"FF979797",
      x"FF888888",
      x"FF717171",
      x"FF565656",
      x"FF353535",
      x"FF111111",
      x"FF000000",
      x"FF000000",
      x"F8000000",
      x"88000000",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"18000000",
      x"C21A1A1A",
      x"FFA7A7A7",
      x"FEE5E5E5",
      x"FFF2F2F2",
      x"FFEEEEEE",
      x"FFE8E8E8",
      x"FFE2E2E2",
      x"FFDCDCDC",
      x"FFD7D7D7",
      x"FFD2D2D2",
      x"FFCECECE",
      x"FFCACACA",
      x"FFC8C8C8",
      x"FFC7C7C7",
      x"FFC6C6C6",
      x"FFC5C5C5",
      x"FFC5C5C5",
      x"FFC6C6C6",
      x"FFC7C7C7",
      x"FFC8C8C8",
      x"FFCACACA",
      x"FFCECECE",
      x"FFD2D2D2",
      x"FFD7D7D7",
      x"FFDCDCDC",
      x"FFE2E2E2",
      x"FFE8E8E8",
      x"FFEEEEEE",
      x"FFF2F2F2",
      x"FEE5E5E5",
      x"FFA8A8A8",
      x"C21E1E1E",
      x"18000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3FA6A6A6",
      x"E8AAAAAA",
      x"FE757575",
      x"FF5A5A5A",
      x"FF4B4B4B",
      x"FF3C3C3C",
      x"FF303030",
      x"FF262626",
      x"FF1E1E1E",
      x"FF181818",
      x"FF111111",
      x"FF0B0B0B",
      x"FF080808",
      x"FF060606",
      x"FF040404",
      x"FF020202",
      x"FF020202",
      x"FF040404",
      x"FF060606",
      x"FF080808",
      x"FF0B0B0B",
      x"FF101010",
      x"FF181818",
      x"FF1E1E1E",
      x"FF262626",
      x"FF303030",
      x"FF3C3C3C",
      x"FF4B4B4B",
      x"FF5A5A5A",
      x"FE757575",
      x"E7A4A4A4",
      x"3FA6A6A6",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01FFFFFF",
      x"5F1E1E1E",
      x"FE040404",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE040404",
      x"5F1B1B1B",
      x"01FFFFFF",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"35000000",
      x"F4000000",
      x"FF000000",
      x"FF020202",
      x"FF050505",
      x"FF080808",
      x"FF0B0B0B",
      x"FF0D0D0D",
      x"FF0F0F0F",
      x"FF111111",
      x"FF151515",
      x"FF181818",
      x"FF1B1B1B",
      x"FF1C1C1C",
      x"FF1D1D1D",
      x"FF1D1D1D",
      x"FF1C1C1C",
      x"FF1B1B1B",
      x"FF181818",
      x"FF151515",
      x"FF111111",
      x"FF0F0F0F",
      x"FF0D0D0D",
      x"FF0B0B0B",
      x"FF080808",
      x"FF050505",
      x"FF020202",
      x"FF000000",
      x"F4000000",
      x"35000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"562F2F2F",
      x"FF3E3E3E",
      x"FF535353",
      x"FF676767",
      x"FF7C7C7C",
      x"FF8C8C8C",
      x"FF9C9C9C",
      x"FFA6A6A6",
      x"FFABABAB",
      x"FFB3B3B3",
      x"FFBBBBBB",
      x"FFC1C1C1",
      x"FFC5C5C5",
      x"FFC7C7C7",
      x"FFCACACA",
      x"FFCACACA",
      x"FFC7C7C7",
      x"FFC5C5C5",
      x"FFC1C1C1",
      x"FFBBBBBB",
      x"FFB3B3B3",
      x"FFABABAB",
      x"FFA6A6A6",
      x"FF9C9C9C",
      x"FF8C8C8C",
      x"FF7B7B7B",
      x"FF676767",
      x"FF535353",
      x"FF404040",
      x"562F2F2F",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"12000000",
      x"D88B8B8B",
      x"FFE9E9E9",
      x"FFF0F0F0",
      x"FFF1F1F1",
      x"FFD7D7D7",
      x"FFB9B9B9",
      x"FF9C9C9C",
      x"FF808080",
      x"FF6B6B6B",
      x"FF595959",
      x"FF474747",
      x"FF3C3C3C",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3C3C3C",
      x"FF484848",
      x"FF5A5A5A",
      x"FF6B6B6B",
      x"FF818181",
      x"FF9D9D9D",
      x"FFB9B9B9",
      x"FFD7D7D7",
      x"FFF1F1F1",
      x"FFF0F0F0",
      x"FFEAEAEA",
      x"D78D8D8D",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"C5000000",
      x"FF1A1A1A",
      x"FF505050",
      x"FF222222",
      x"FF000000",
      x"FF010101",
      x"FF030303",
      x"FF050505",
      x"FF060606",
      x"FF070707",
      x"FF090909",
      x"FF0A0A0A",
      x"FF0A0A0A",
      x"FF0A0A0A",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0B0B0B",
      x"FF0A0A0A",
      x"FF0A0A0A",
      x"FF0A0A0A",
      x"FF090909",
      x"FF080808",
      x"FF070707",
      x"FF050505",
      x"FF040404",
      x"FF020202",
      x"FF000000",
      x"FF000000",
      x"FF232323",
      x"FF4E4E4E",
      x"FF191919",
      x"B5000000",
      x"06000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"5F000000",
      x"F2111111",
      x"FF282828",
      x"FF3B3B3B",
      x"FF4B4B4B",
      x"FF565656",
      x"FF606060",
      x"FF6E6E6E",
      x"FF797979",
      x"FF808080",
      x"FF888888",
      x"FF909090",
      x"FF969696",
      x"FF989898",
      x"FF9B9B9B",
      x"FF9D9D9D",
      x"FF9F9F9F",
      x"FF9F9F9F",
      x"FF9C9C9C",
      x"FF999999",
      x"FF979797",
      x"FF939393",
      x"FF8B8B8B",
      x"FF838383",
      x"FF7B7B7B",
      x"FF727272",
      x"FF656565",
      x"FF595959",
      x"FF4F4F4F",
      x"FF424242",
      x"FF2F2F2F",
      x"FF181818",
      x"E1030303",
      x"32000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0B8B8B8B",
      x"99ACACAC",
      x"FDCBCBCB",
      x"FFDDDDDD",
      x"FFE8E8E8",
      x"FFEDEDED",
      x"FFF1F1F1",
      x"FFF3F3F3",
      x"FFEAEAEA",
      x"FFDADADA",
      x"FFCDCDCD",
      x"FFC0C0C0",
      x"FFB3B3B3",
      x"FFA9A9A9",
      x"FFA3A3A3",
      x"FFA1A1A1",
      x"FF9C9C9C",
      x"FF979797",
      x"FF9C9C9C",
      x"FF9F9F9F",
      x"FFA1A1A1",
      x"FFA9A9A9",
      x"FFAEAEAE",
      x"FFBBBBBB",
      x"FFC9C9C9",
      x"FFD6D6D6",
      x"FFE5E5E5",
      x"FFF4F4F4",
      x"FFF2F2F2",
      x"FFEFEFEF",
      x"FFEAEAEA",
      x"FFE1E1E1",
      x"FFD2D2D2",
      x"EBB4B4B4",
      x"475A5A5A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"29252525",
      x"E0737373",
      x"FEB5B5B5",
      x"FF878787",
      x"FF595959",
      x"FF353535",
      x"FF191919",
      x"FF030303",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF010101",
      x"FF0F0F0F",
      x"FF2C2C2C",
      x"FF4B4B4B",
      x"FF777777",
      x"FFACACAC",
      x"F9A7A7A7",
      x"80323232",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3B000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"AF000000",
      x"10000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"25000000",
      x"D9000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"A2000000",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"04000000",
      x"5D000000",
      x"D6000000",
      x"E9000000",
      x"F1000000",
      x"F5000000",
      x"F8000000",
      x"FA000000",
      x"FC000000",
      x"FE000000",
      x"FF000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"FF000000",
      x"FE000000",
      x"FC000000",
      x"FA000000",
      x"F8000000",
      x"F5000000",
      x"F1000000",
      x"E9000000",
      x"D2000000",
      x"46000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"2A000000",
      x"45000000",
      x"56000000",
      x"68000000",
      x"7A000000",
      x"87000000",
      x"95000000",
      x"A2000000",
      x"A9000000",
      x"AF000000",
      x"B6000000",
      x"BD000000",
      x"C1000000",
      x"C4000000",
      x"C6000000",
      x"C9000000",
      x"CA000000",
      x"C6000000",
      x"C4000000",
      x"C1000000",
      x"BD000000",
      x"B6000000",
      x"AF000000",
      x"A9000000",
      x"A2000000",
      x"95000000",
      x"87000000",
      x"7A000000",
      x"68000000",
      x"56000000",
      x"45000000",
      x"2C000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"05000000",
      x"08000000",
      x"0A000000",
      x"0C000000",
      x"0E000000",
      x"10000000",
      x"13000000",
      x"17000000",
      x"19000000",
      x"1A000000",
      x"1B000000",
      x"1D000000",
      x"1D000000",
      x"1C000000",
      x"1A000000",
      x"19000000",
      x"17000000",
      x"13000000",
      x"10000000",
      x"0E000000",
      x"0C000000",
      x"0A000000",
      x"08000000",
      x"05000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
