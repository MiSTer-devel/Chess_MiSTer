library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_white_pawn_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_white_pawn_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"29000000",
      x"32000000",
      x"21000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"5F000000",
      x"C9000000",
      x"DA000000",
      x"DF000000",
      x"D6000000",
      x"AA000000",
      x"25000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"15000000",
      x"9D000000",
      x"FB000000",
      x"FE090909",
      x"FF161616",
      x"FF1C1C1C",
      x"FE111111",
      x"FE050505",
      x"FF000000",
      x"62000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"04000000",
      x"9A000000",
      x"FA000000",
      x"FF313131",
      x"FF8D8D8D",
      x"FFBBBBBB",
      x"FFC8C8C8",
      x"FFB0B0B0",
      x"FF6D6D6D",
      x"FE0C0C0C",
      x"F1000000",
      x"62000000",
      x"04000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"66000000",
      x"FA000000",
      x"FF333333",
      x"FFCDCDCD",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF969696",
      x"FF000000",
      x"C7000000",
      x"1E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"06000000",
      x"C8000000",
      x"FE090909",
      x"FF8B8B8B",
      x"FFFAFAFA",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF464646",
      x"FE000000",
      x"43000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"27000000",
      x"D9000000",
      x"FF161616",
      x"FFBCBCBC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFB1B1B1",
      x"FF000000",
      x"7A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"30000000",
      x"DF000000",
      x"FF1C1C1C",
      x"FFC6C6C6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFC3C3C3",
      x"FF000000",
      x"8E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1E000000",
      x"D4000000",
      x"FE121212",
      x"FFB1B1B1",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FF9D9D9D",
      x"FF000000",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"AC000000",
      x"FF040404",
      x"FF6B6B6B",
      x"FFF3F3F3",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFE2E2E2",
      x"FF262626",
      x"EF000000",
      x"32000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1D000000",
      x"C7000000",
      x"FF000000",
      x"FF0D0D0D",
      x"FFC5C5C5",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFBFBFB",
      x"FF515151",
      x"FF000000",
      x"FA000000",
      x"6B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"A5000000",
      x"FC000000",
      x"FF1A1A1A",
      x"FF8B8B8B",
      x"FFF6F6F6",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFECECEC",
      x"FF525252",
      x"FE0D0D0D",
      x"FF000000",
      x"6C000000",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"84000000",
      x"F6000000",
      x"FF363636",
      x"FFBBBBBB",
      x"FFFCFCFC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF5F5F5",
      x"FF8C8C8C",
      x"FE0E0E0E",
      x"ED000000",
      x"53000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"42000000",
      x"F6000000",
      x"FE252525",
      x"FFC7C7C7",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF7F7F7",
      x"FF747474",
      x"FE000000",
      x"B4000000",
      x"15000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"C0000000",
      x"FF050505",
      x"FF787878",
      x"FFF7F7F7",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF232323",
      x"F6000000",
      x"3E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2E000000",
      x"DD000000",
      x"FF171717",
      x"FFBCBCBC",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFA5A5A5",
      x"FE030303",
      x"89000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"50000000",
      x"EE000000",
      x"FF2D2D2D",
      x"FFE6E6E6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFD3D3D3",
      x"FF1D1D1D",
      x"D6000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"5D000000",
      x"F3000000",
      x"FF373737",
      x"FFF8F8F8",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFDDDDDD",
      x"FF2F2F2F",
      x"FB000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"5E000000",
      x"F3000000",
      x"FF373737",
      x"FFF9F9F9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFDDDDDD",
      x"FF2F2F2F",
      x"FA000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"50000000",
      x"EF000000",
      x"FF2D2D2D",
      x"FFE7E7E7",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFD3D3D3",
      x"FF1D1D1D",
      x"D6000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"30000000",
      x"DF000000",
      x"FE171717",
      x"FFBCBCBC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFACACAC",
      x"FF000000",
      x"8F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"B7000000",
      x"FE050505",
      x"FF787878",
      x"FFF7F7F7",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF1F1F1",
      x"FF313131",
      x"F2000000",
      x"40000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"36000000",
      x"FF000000",
      x"FE1C1C1C",
      x"FFD3D3D3",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FF6C6C6C",
      x"FF010101",
      x"B7000000",
      x"14000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"85000000",
      x"FB000000",
      x"FF232323",
      x"FFD7D7D7",
      x"FFFBFBFB",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF5F5F5",
      x"FF959595",
      x"FF0D0D0D",
      x"EE000000",
      x"56000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"60000000",
      x"ED000000",
      x"FF000000",
      x"FF262626",
      x"FFB1B1B1",
      x"FFFCFCFC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFCFCFC",
      x"FF858585",
      x"FF161616",
      x"FF000000",
      x"DF000000",
      x"3D000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"9A000000",
      x"ED000000",
      x"FD000000",
      x"FF191919",
      x"FF8C8C8C",
      x"FFDEDEDE",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FFC7C7C7",
      x"FF626262",
      x"FF080808",
      x"FC000000",
      x"DB000000",
      x"48000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"14000000",
      x"9B000000",
      x"FB000000",
      x"FE131313",
      x"FF727272",
      x"FFF1F1F1",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD2D2D2",
      x"FF3B3B3B",
      x"FE080808",
      x"FF000000",
      x"5D000000",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0B000000",
      x"99000000",
      x"F7000000",
      x"FF2F2F2F",
      x"FFA8A8A8",
      x"FFF5F5F5",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFEFEFEF",
      x"FF7C7C7C",
      x"FE0C0C0C",
      x"F0000000",
      x"62000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"95000000",
      x"FA000000",
      x"FF2F2F2F",
      x"FFCACACA",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF5F5F5",
      x"FF8F8F8F",
      x"FF000000",
      x"E3000000",
      x"2F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"55000000",
      x"EE000000",
      x"FE141414",
      x"FFABABAB",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF7B7B7B",
      x"FE060606",
      x"CC000000",
      x"10000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"17000000",
      x"B9000000",
      x"FD000000",
      x"FF7B7B7B",
      x"FFF6F6F6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFECECEC",
      x"FF4D4D4D",
      x"FF020202",
      x"93000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"58000000",
      x"F9000000",
      x"FE3B3B3B",
      x"FFF4F4F4",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFB0B0B0",
      x"FE131313",
      x"E7000000",
      x"42000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"E0000000",
      x"FF090909",
      x"FFC3C3C3",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF8F8F8",
      x"FF4A4A4A",
      x"FA000000",
      x"8D000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"67000000",
      x"FF010101",
      x"FE4D4D4D",
      x"FFEBEBEB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFC9C9C9",
      x"FF030303",
      x"CB000000",
      x"1E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0A000000",
      x"C2000000",
      x"FF090909",
      x"FF8E8E8E",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FF4E4E4E",
      x"FA000000",
      x"41000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"35000000",
      x"E1000000",
      x"FF181818",
      x"FFC0C0C0",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFB7B7B7",
      x"FF030303",
      x"99000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"5A000000",
      x"F1000000",
      x"FF323232",
      x"FFEFEFEF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD9D9D9",
      x"FF252525",
      x"E8000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"06000000",
      x"7C000000",
      x"F8000000",
      x"FF5B5B5B",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFECECEC",
      x"FF4A4A4A",
      x"FF000000",
      x"28000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0B000000",
      x"99000000",
      x"FD000000",
      x"FF969696",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF626262",
      x"FF020202",
      x"65000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"AD000000",
      x"FF000000",
      x"FFC5C5C5",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF8F8F8",
      x"FF797979",
      x"FF050505",
      x"95000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"16000000",
      x"BC000000",
      x"FE000000",
      x"FFE9E9E9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFAFAFA",
      x"FF8B8B8B",
      x"FF080808",
      x"B8000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1A000000",
      x"C4000000",
      x"FF000000",
      x"FFC0C0C0",
      x"FFC4C4C4",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC2C2C2",
      x"FF717171",
      x"FE070707",
      x"C3000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1E000000",
      x"CA000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C8000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"11000000",
      x"78000000",
      x"96000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"95000000",
      x"74000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
