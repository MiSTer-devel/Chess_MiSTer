library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_tile_1 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_tile_1 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"FFF2A34A",
      x"FFF2A14A",
      x"FFF3A550",
      x"FFEC953B",
      x"FFE9903A",
      x"FFEA943D",
      x"FFEE9D4C",
      x"FFEC9D4F",
      x"FFE99748",
      x"FFE58C38",
      x"FFE89438",
      x"FFF4A638",
      x"FFF9AE3A",
      x"FFFAAB37",
      x"FFFCB03F",
      x"FFFAB348",
      x"FFF89E29",
      x"FFFA9F28",
      x"FFF7A030",
      x"FFF79E2F",
      x"FFF69A24",
      x"FFFAA830",
      x"FFFDAC2C",
      x"FFFAAD41",
      x"FFFBA937",
      x"FFF8A12D",
      x"FFFDB954",
      x"FFFDBD51",
      x"FFFDB33B",
      x"FFF8A525",
      x"FFE88C1F",
      x"FFD67014",
      x"FFD7731C",
      x"FFE08124",
      x"FFDF8023",
      x"FFDF8524",
      x"FFD97922",
      x"FFDB7B1E",
      x"FFDC7E22",
      x"FFDC8426",
      x"FFD37C23",
      x"FFD37A20",
      x"FFD68224",
      x"FFD78624",
      x"FFD27D21",
      x"FFD67D20",
      x"FFDC8A28",
      x"FFE09230",
      x"FFD78B30",
      x"FFD48C34",
      x"FFCC8430",
      x"FFD08633",
      x"FFD78E40",
      x"FFDD8F4A",
      x"FFDC934B",
      x"FFD98E41",
      x"FFD38634",
      x"FFD17E29",
      x"FFCE7723",
      x"FFCD741E",
      x"FFF0A24B",
      x"FFF1A14A",
      x"FFF3A34E",
      x"FFED9741",
      x"FFEC9742",
      x"FFE98E36",
      x"FFEC9A49",
      x"FFEDA35B",
      x"FFE99748",
      x"FFE99445",
      x"FFE68F36",
      x"FFEEA13C",
      x"FFF9B140",
      x"FFFAAD39",
      x"FFFBAC38",
      x"FFFCB752",
      x"FFFAAB3E",
      x"FFFBA22A",
      x"FFF9A129",
      x"FFF6A136",
      x"FFF69C25",
      x"FFF8A129",
      x"FFFBAE37",
      x"FFFBB03F",
      x"FFFBA737",
      x"FFFBA936",
      x"FFFBB148",
      x"FFFCB951",
      x"FFFDBC51",
      x"FFF8A123",
      x"FFEB8E1C",
      x"FFD77213",
      x"FFD57019",
      x"FFDF7D20",
      x"FFE08223",
      x"FFDF7F21",
      x"FFD7751E",
      x"FFDC7C20",
      x"FFDC7A1D",
      x"FFDD8326",
      x"FFD57D23",
      x"FFD07720",
      x"FFD47E21",
      x"FFD78223",
      x"FFD47E21",
      x"FFD98123",
      x"FFDA8525",
      x"FFDF9333",
      x"FFD88C2E",
      x"FFD58D35",
      x"FFCC812B",
      x"FFCA7C2C",
      x"FFD48C3A",
      x"FFD98F48",
      x"FFDA9148",
      x"FFDA9044",
      x"FFD48736",
      x"FFD0812C",
      x"FFCC7824",
      x"FFCD721E",
      x"FFF1A550",
      x"FFF0A04A",
      x"FFF09E49",
      x"FFEF9D49",
      x"FFED9945",
      x"FFE88D39",
      x"FFEE9C4B",
      x"FFEDA25A",
      x"FFEC9D51",
      x"FFE89343",
      x"FFE8933F",
      x"FFEA993D",
      x"FFF6AF45",
      x"FFFBAE3B",
      x"FFFBAC38",
      x"FFFCB247",
      x"FFFBAF42",
      x"FFF99D26",
      x"FFFBAB3B",
      x"FFF8A436",
      x"FFF59A25",
      x"FFF69923",
      x"FFFAA82F",
      x"FFFBAF38",
      x"FFFAA736",
      x"FFFAA939",
      x"FFFAAB40",
      x"FFFBB045",
      x"FFFDBB55",
      x"FFF9AA32",
      x"FFEC8D1C",
      x"FFDA7716",
      x"FFD46B17",
      x"FFDD7B20",
      x"FFE18526",
      x"FFDD7D1F",
      x"FFD87921",
      x"FFDA771C",
      x"FFDA771B",
      x"FFDC8123",
      x"FFD57E25",
      x"FFD0751D",
      x"FFD27B1F",
      x"FFD88424",
      x"FFD58125",
      x"FFD77D20",
      x"FFDA8525",
      x"FFE29632",
      x"FFDA8E31",
      x"FFD38A31",
      x"FFCF862E",
      x"FFC87B29",
      x"FFD48A37",
      x"FFD68D44",
      x"FFDB9147",
      x"FFD98F44",
      x"FFD58735",
      x"FFD1822E",
      x"FFCC7422",
      x"FFCE731E",
      x"FFF1A14D",
      x"FFF19F4A",
      x"FFF19F4D",
      x"FFEF9C4C",
      x"FFED9441",
      x"FFE98F3C",
      x"FFED9846",
      x"FFEDA157",
      x"FFEC9C51",
      x"FFE7903D",
      x"FFE38C3C",
      x"FFE7953C",
      x"FFEFA540",
      x"FFF9B444",
      x"FFFBAD3C",
      x"FFFAAC3A",
      x"FFFCB146",
      x"FFFBA12A",
      x"FFFBAE3F",
      x"FFFAAC41",
      x"FFF59E30",
      x"FFF38F1B",
      x"FFF89C21",
      x"FFFAAF3B",
      x"FFFAAA38",
      x"FFF9A22D",
      x"FFF9A93A",
      x"FFF9A42F",
      x"FFFAAE3A",
      x"FFF9B13D",
      x"FFEC9021",
      x"FFDD7915",
      x"FFD16711",
      x"FFDB7A20",
      x"FFDF8425",
      x"FFDC781B",
      x"FFDA7B22",
      x"FFDD7D20",
      x"FFDA791D",
      x"FFDF8224",
      x"FFD57D23",
      x"FFD17820",
      x"FFD27C20",
      x"FFD88322",
      x"FFD88324",
      x"FFD57E21",
      x"FFD88122",
      x"FFE39532",
      x"FFD98E31",
      x"FFD48B30",
      x"FFD18931",
      x"FFCD7F2B",
      x"FFD28631",
      x"FFD68F42",
      x"FFD99148",
      x"FFDA9046",
      x"FFD68537",
      x"FFD48430",
      x"FFCC731F",
      x"FFCB731E",
      x"FFED9941",
      x"FFF1A34E",
      x"FFF2A655",
      x"FFF2A353",
      x"FFEE9743",
      x"FFEC9646",
      x"FFEE9741",
      x"FFEFA358",
      x"FFED9E51",
      x"FFEA933C",
      x"FFE99441",
      x"FFE79139",
      x"FFEEA347",
      x"FFF7B145",
      x"FFFBB042",
      x"FFFBAB39",
      x"FFFCB44C",
      x"FFFAA534",
      x"FFFBAB38",
      x"FFFAA939",
      x"FFF7A63B",
      x"FFF28D1C",
      x"FFF6951F",
      x"FFF9A42D",
      x"FFFAAA35",
      x"FFF7A12D",
      x"FFF9A430",
      x"FFF9A027",
      x"FFF6A328",
      x"FFFAB03B",
      x"FFEC8E1C",
      x"FFE3851D",
      x"FFD06411",
      x"FFD8721A",
      x"FFDE7F22",
      x"FFDC791D",
      x"FFDA7C21",
      x"FFDE8023",
      x"FFDA781D",
      x"FFDC7F21",
      x"FFD87F24",
      x"FFD27920",
      x"FFD0791E",
      x"FFD88324",
      x"FFD88123",
      x"FFD88022",
      x"FFD87F21",
      x"FFE39735",
      x"FFDB9031",
      x"FFD5892E",
      x"FFD28931",
      x"FFCC802C",
      x"FFCF812F",
      x"FFD89143",
      x"FFD78F44",
      x"FFD99246",
      x"FFD48535",
      x"FFD78B35",
      x"FFCB721F",
      x"FFCC721E",
      x"FFEB9842",
      x"FFF2A24D",
      x"FFF09F4B",
      x"FFF2A453",
      x"FFEE9944",
      x"FFEE9641",
      x"FFEC953F",
      x"FFF1A658",
      x"FFEC9E50",
      x"FFE69247",
      x"FFE79345",
      x"FFE78E3C",
      x"FFE99A42",
      x"FFF4AB40",
      x"FFFAB146",
      x"FFFBB143",
      x"FFFCB854",
      x"FFFAAD41",
      x"FFFBA933",
      x"FFFBA936",
      x"FFFAB04A",
      x"FFF39427",
      x"FFF5921B",
      x"FFF89D25",
      x"FFF9A733",
      x"FFF8A22D",
      x"FFF8A32D",
      x"FFF8A42D",
      x"FFF8A327",
      x"FFF9A82A",
      x"FFEE9422",
      x"FFE5891F",
      x"FFD16A12",
      x"FFD66D16",
      x"FFDD7D1F",
      x"FFDA7319",
      x"FFDC7E21",
      x"FFDB781F",
      x"FFD8751B",
      x"FFDC7E22",
      x"FFD87D22",
      x"FFCF7920",
      x"FFD37B1F",
      x"FFD68123",
      x"FFD78224",
      x"FFD67E21",
      x"FFD67E20",
      x"FFE29330",
      x"FFDB8F30",
      x"FFD3862A",
      x"FFD2872D",
      x"FFCA7E27",
      x"FFCC7F2B",
      x"FFD58E40",
      x"FFD79046",
      x"FFD9944A",
      x"FFD88C3F",
      x"FFD48834",
      x"FFCE7821",
      x"FFCC721E",
      x"FFE7923E",
      x"FFF1A350",
      x"FFF09F4B",
      x"FFF19F4A",
      x"FFEC9945",
      x"FFEC953E",
      x"FFEA933D",
      x"FFF1A251",
      x"FFEEA154",
      x"FFE59043",
      x"FFE69448",
      x"FFE58B38",
      x"FFE99946",
      x"FFF0A647",
      x"FFFAB349",
      x"FFFBB042",
      x"FFFCB54D",
      x"FFFBB451",
      x"FFFBAB37",
      x"FFFCA329",
      x"FFFBAD41",
      x"FFF49D34",
      x"FFF48E1C",
      x"FFF6981E",
      x"FFF69F2B",
      x"FFF69C26",
      x"FFF9A634",
      x"FFF9A22A",
      x"FFFAA528",
      x"FFF89F20",
      x"FFF29824",
      x"FFE68519",
      x"FFD46B13",
      x"FFD6731A",
      x"FFDF8022",
      x"FFD9771D",
      x"FFDE8123",
      x"FFD97820",
      x"FFD9751A",
      x"FFDC7F23",
      x"FFD98023",
      x"FFD0771F",
      x"FFD17A20",
      x"FFD58023",
      x"FFD88222",
      x"FFD67F20",
      x"FFD87F20",
      x"FFE29130",
      x"FFDD9032",
      x"FFD78F35",
      x"FFD28930",
      x"FFCE822A",
      x"FFCA7E2B",
      x"FFD38837",
      x"FFD78F45",
      x"FFD89449",
      x"FFD88F41",
      x"FFD38533",
      x"FFCF7923",
      x"FFCD7420",
      x"FFE89137",
      x"FFED9A45",
      x"FFF2A14C",
      x"FFEF9C49",
      x"FFED9741",
      x"FFEB9039",
      x"FFEA913C",
      x"FFED9B46",
      x"FFEEA254",
      x"FFE79648",
      x"FFE89445",
      x"FFE78E41",
      x"FFE7913F",
      x"FFEDA44E",
      x"FFF6AD45",
      x"FFFBB44C",
      x"FFFCB448",
      x"FFFCBD61",
      x"FFFBAF45",
      x"FFFAA229",
      x"FFFAA738",
      x"FFF6A134",
      x"FFF59422",
      x"FFF69B23",
      x"FFF79F28",
      x"FFF59826",
      x"FFF8A533",
      x"FFF89E26",
      x"FFF9A329",
      x"FFF8A122",
      x"FFF08F19",
      x"FFE68719",
      x"FFD4680E",
      x"FFD66F18",
      x"FFDD7C20",
      x"FFD9721A",
      x"FFDE8022",
      x"FFD77621",
      x"FFDC7A1F",
      x"FFDC7D21",
      x"FFD87F24",
      x"FFD2781F",
      x"FFD1791F",
      x"FFD57F23",
      x"FFD88424",
      x"FFD47A1D",
      x"FFD98122",
      x"FFDF8E2B",
      x"FFE09434",
      x"FFD68C32",
      x"FFD38C34",
      x"FFCE8530",
      x"FFCC8430",
      x"FFD28534",
      x"FFD99245",
      x"FFD99347",
      x"FFD78F40",
      x"FFD28331",
      x"FFD27E28",
      x"FFCC741F",
      x"FFE9953B",
      x"FFEB953D",
      x"FFF09E46",
      x"FFEE9D49",
      x"FFED9741",
      x"FFEC943E",
      x"FFEB9441",
      x"FFEA943F",
      x"FFF0A353",
      x"FFEA9A4C",
      x"FFE99344",
      x"FFE89447",
      x"FFE68E3E",
      x"FFECA150",
      x"FFF1A641",
      x"FFFBB64F",
      x"FFFBB243",
      x"FFFCBB5C",
      x"FFFAA83A",
      x"FFFBAC3B",
      x"FFF9A42E",
      x"FFF79D2C",
      x"FFF39423",
      x"FFF59D29",
      x"FFF39A26",
      x"FFF39421",
      x"FFF69F29",
      x"FFF7A029",
      x"FFF89F25",
      x"FFF8A123",
      x"FFF28C13",
      x"FFE9881B",
      x"FFD5680E",
      x"FFD46C15",
      x"FFDB771B",
      x"FFD9741B",
      x"FFDF7F20",
      x"FFD6741C",
      x"FFDB7A1F",
      x"FFDC7C1F",
      x"FFDB8023",
      x"FFD57C22",
      x"FFD17A1F",
      x"FFD47E22",
      x"FFD78425",
      x"FFD67D1F",
      x"FFDA8423",
      x"FFDE8824",
      x"FFE19836",
      x"FFD78B30",
      x"FFD68F36",
      x"FFCF8734",
      x"FFD08834",
      x"FFD08535",
      x"FFD99143",
      x"FFDB9548",
      x"FFDA9242",
      x"FFD18130",
      x"FFCF7D26",
      x"FFCE7521",
      x"FFE8943E",
      x"FFE88E35",
      x"FFED9840",
      x"FFF09B46",
      x"FFF19E4A",
      x"FFEA8E38",
      x"FFEC933E",
      x"FFE8903A",
      x"FFF1A24E",
      x"FFEEA254",
      x"FFE99548",
      x"FFE89549",
      x"FFE79141",
      x"FFEB994A",
      x"FFEEA44B",
      x"FFF7B24A",
      x"FFFCB54A",
      x"FFFCBB56",
      x"FFFAAC3D",
      x"FFFDB549",
      x"FFFBA530",
      x"FFF79B26",
      x"FFF3901E",
      x"FFF59E2E",
      x"FFF49D2C",
      x"FFEF8F20",
      x"FFF38E17",
      x"FFF8A02A",
      x"FFF3951F",
      x"FFF79F28",
      x"FFF38D14",
      x"FFED8A19",
      x"FFD66C0E",
      x"FFD36A13",
      x"FFD87319",
      x"FFDB7A1D",
      x"FFDE7C1F",
      x"FFD4731C",
      x"FFDA791E",
      x"FFD8771C",
      x"FFDC8124",
      x"FFD37A21",
      x"FFD0781D",
      x"FFD57D20",
      x"FFD47E22",
      x"FFD78022",
      x"FFDB8120",
      x"FFDB8321",
      x"FFE29735",
      x"FFD88E32",
      x"FFD48D34",
      x"FFCE8634",
      x"FFD08934",
      x"FFCC802E",
      x"FFD89040",
      x"FFDC9549",
      x"FFD89041",
      x"FFD28332",
      x"FFCF7E27",
      x"FFCE7722",
      x"FFEB973F",
      x"FFE4882F",
      x"FFEA953F",
      x"FFEE9B46",
      x"FFF1A24E",
      x"FFEB943D",
      x"FFE8913C",
      x"FFE88F3A",
      x"FFF19F48",
      x"FFF0A353",
      x"FFEB994B",
      x"FFEA9B51",
      x"FFE58F41",
      x"FFEA994A",
      x"FFEEA24D",
      x"FFF6B14F",
      x"FFFBB755",
      x"FFFCBC5C",
      x"FFFAAF46",
      x"FFFCB752",
      x"FFFBAA35",
      x"FFF89F29",
      x"FFF6941D",
      x"FFF59625",
      x"FFF29D2E",
      x"FFF09527",
      x"FFF08410",
      x"FFF4921C",
      x"FFF08F1E",
      x"FFF79D25",
      x"FFF6961B",
      x"FFEC8514",
      x"FFD86D0F",
      x"FFD46A13",
      x"FFD66F16",
      x"FFDB771B",
      x"FFDB771C",
      x"FFD6761D",
      x"FFD9771C",
      x"FFD77419",
      x"FFDE8427",
      x"FFD37C22",
      x"FFD2781F",
      x"FFD27A1F",
      x"FFD58226",
      x"FFD27B21",
      x"FFD77B1D",
      x"FFDA8120",
      x"FFE29937",
      x"FFDA8F35",
      x"FFD58D36",
      x"FFD18C3A",
      x"FFCE8633",
      x"FFC98030",
      x"FFD4893B",
      x"FFDC9649",
      x"FFD88F3F",
      x"FFD58835",
      x"FFD2832C",
      x"FFCB721D",
      x"FFEB973E",
      x"FFE78C32",
      x"FFEB953D",
      x"FFED9942",
      x"FFF2A14B",
      x"FFED923A",
      x"FFEB913B",
      x"FFE78D3A",
      x"FFF09D45",
      x"FFF1A351",
      x"FFEB9B4B",
      x"FFE79245",
      x"FFE59244",
      x"FFE99344",
      x"FFEC9F4C",
      x"FFF1A950",
      x"FFF9B651",
      x"FFFCBD61",
      x"FFFBB54B",
      x"FFFDB64D",
      x"FFFCB142",
      x"FFF9A42E",
      x"FFF5951F",
      x"FFF6921D",
      x"FFF19D31",
      x"FFEF9829",
      x"FFF08514",
      x"FFE87C10",
      x"FFF49821",
      x"FFF4971E",
      x"FFF79A1F",
      x"FFE97C0C",
      x"FFDF730E",
      x"FFD26913",
      x"FFD36913",
      x"FFDB771B",
      x"FFDA761A",
      x"FFD97A1F",
      x"FFDB771C",
      x"FFD77117",
      x"FFDC8225",
      x"FFD37A20",
      x"FFD2791F",
      x"FFD57E22",
      x"FFD68226",
      x"FFD27E21",
      x"FFD97C1B",
      x"FFDA7E1D",
      x"FFE49936",
      x"FFD98E33",
      x"FFD58E37",
      x"FFD18B38",
      x"FFCB8532",
      x"FFCB8232",
      x"FFD08535",
      x"FFDC9447",
      x"FFD78E3E",
      x"FFD68632",
      x"FFD2832D",
      x"FFCF7B22",
      x"FFEA9338",
      x"FFE5872C",
      x"FFEA9238",
      x"FFEB933A",
      x"FFF09A42",
      x"FFF09940",
      x"FFEC9139",
      x"FFEA9442",
      x"FFEC9741",
      x"FFF2A454",
      x"FFEEA153",
      x"FFE79548",
      x"FFE99447",
      x"FFE89545",
      x"FFEB9C4B",
      x"FFECA34D",
      x"FFF6B04F",
      x"FFF9B653",
      x"FFFCB64B",
      x"FFFBB042",
      x"FFFDB64E",
      x"FFF8A531",
      x"FFF79B1F",
      x"FFF6901A",
      x"FFF19727",
      x"FFEF972C",
      x"FFEC8818",
      x"FFE87608",
      x"FFF38C16",
      x"FFF89C21",
      x"FFF79C1F",
      x"FFED8512",
      x"FFE17811",
      x"FFD1630D",
      x"FFD46E16",
      x"FFDD7B1D",
      x"FFDA751A",
      x"FFDC7D22",
      x"FFD9781E",
      x"FFD87219",
      x"FFDC7F22",
      x"FFD37B21",
      x"FFD1761D",
      x"FFD27B21",
      x"FFD07B23",
      x"FFD37D21",
      x"FFD77D1E",
      x"FFDA7F1F",
      x"FFE39734",
      x"FFDA8E34",
      x"FFD89039",
      x"FFD28A38",
      x"FFD18933",
      x"FFD08836",
      x"FFD08533",
      x"FFDA9348",
      x"FFD99040",
      x"FFD78A38",
      x"FFD28530",
      x"FFD08028",
      x"FFE99135",
      x"FFE5882C",
      x"FFEB9134",
      x"FFEB9036",
      x"FFED9840",
      x"FFF29E47",
      x"FFED933C",
      x"FFEC953D",
      x"FFED953C",
      x"FFF2A24E",
      x"FFF1A456",
      x"FFEB9D50",
      x"FFE89549",
      x"FFE79444",
      x"FFEC9B49",
      x"FFEB9C4B",
      x"FFF4AD53",
      x"FFF9B654",
      x"FFFBB54A",
      x"FFFBB042",
      x"FFFDBD5A",
      x"FFF9AC40",
      x"FFFAA123",
      x"FFF5901A",
      x"FFF2911E",
      x"FFEE9527",
      x"FFEC8C20",
      x"FFEF820E",
      x"FFF3860D",
      x"FFF5931D",
      x"FFF5961C",
      x"FFEF8711",
      x"FFE58215",
      x"FFD3630C",
      x"FFD57116",
      x"FFDA781D",
      x"FFD97118",
      x"FFDC7E20",
      x"FFDA791D",
      x"FFD87117",
      x"FFD87D21",
      x"FFD3771F",
      x"FFD0761E",
      x"FFD17A21",
      x"FFD47E23",
      x"FFD37E22",
      x"FFD77C1E",
      x"FFDC801E",
      x"FFE39532",
      x"FFDC9135",
      x"FFD89039",
      x"FFD38C38",
      x"FFD48E39",
      x"FFD08734",
      x"FFCD8334",
      x"FFD88F3F",
      x"FFD99042",
      x"FFDA8D39",
      x"FFD3852F",
      x"FFD3852C",
      x"FFE88C31",
      x"FFE88C32",
      x"FFEA9133",
      x"FFEC9237",
      x"FFEA943C",
      x"FFF09C45",
      x"FFEE943B",
      x"FFEC943E",
      x"FFEC9139",
      x"FFF3A14A",
      x"FFF3A95A",
      x"FFEEA357",
      x"FFE79547",
      x"FFE79243",
      x"FFEA9747",
      x"FFEB9B49",
      x"FFEFA754",
      x"FFF7B354",
      x"FFFBBA5B",
      x"FFFBAB36",
      x"FFFDBC57",
      x"FFFCBA56",
      x"FFF9A228",
      x"FFF48E18",
      x"FFF48D17",
      x"FFED8F24",
      x"FFEC8D21",
      x"FFEE8717",
      x"FFF3870D",
      x"FFF39018",
      x"FFF69418",
      x"FFF18F16",
      x"FFE88216",
      x"FFD76F11",
      x"FFD56D14",
      x"FFD97419",
      x"FFD87319",
      x"FFDE8021",
      x"FFDB791D",
      x"FFD87317",
      x"FFDB7D20",
      x"FFCF741E",
      x"FFCF761E",
      x"FFD07922",
      x"FFD47F23",
      x"FFD47F21",
      x"FFD87D1E",
      x"FFDC811F",
      x"FFE08E2C",
      x"FFDB9032",
      x"FFD8903A",
      x"FFD48B38",
      x"FFD4903B",
      x"FFD18937",
      x"FFCE8634",
      x"FFD58C3C",
      x"FFD78D3E",
      x"FFDA8D3B",
      x"FFD5862E",
      x"FFD18126",
      x"FFEA933A",
      x"FFEB9337",
      x"FFE98C2E",
      x"FFEC9439",
      x"FFE88E34",
      x"FFED9640",
      x"FFF09C44",
      x"FFED9238",
      x"FFEA9039",
      x"FFF2A048",
      x"FFF3A450",
      x"FFEFA253",
      x"FFE79648",
      x"FFE79143",
      x"FFE99547",
      x"FFED9E4B",
      x"FFEDA14E",
      x"FFF5B258",
      x"FFF9B550",
      x"FFFBB146",
      x"FFFCB043",
      x"FFFDC161",
      x"FFFBAB39",
      x"FFF58F17",
      x"FFF38B14",
      x"FFF19120",
      x"FFED9329",
      x"FFEA8115",
      x"FFF18A14",
      x"FFF49219",
      x"FFF5951D",
      x"FFF08D17",
      x"FFE98213",
      x"FFD96F0F",
      x"FFD46B11",
      x"FFD87218",
      x"FFD77218",
      x"FFDE7F1F",
      x"FFD77419",
      x"FFD97318",
      x"FFDB7B1E",
      x"FFCF721D",
      x"FFCF741D",
      x"FFD07720",
      x"FFD37D22",
      x"FFD58329",
      x"FFD87D1E",
      x"FFDF8521",
      x"FFE4922D",
      x"FFDB9135",
      x"FFD88F39",
      x"FFD58C3A",
      x"FFD48F3A",
      x"FFD18B37",
      x"FFCF8735",
      x"FFD38836",
      x"FFDA9345",
      x"FFD98A38",
      x"FFD78832",
      x"FFD17E25",
      x"FFE89038",
      x"FFEA9138",
      x"FFE5862A",
      x"FFEB9235",
      x"FFEA9236",
      x"FFEA913A",
      x"FFEC933B",
      x"FFEE963B",
      x"FFED963E",
      x"FFF29E46",
      x"FFF4A652",
      x"FFF2A452",
      x"FFE79443",
      x"FFE79346",
      x"FFE58F41",
      x"FFED9D4D",
      x"FFEB9F4C",
      x"FFF0AA57",
      x"FFF8B451",
      x"FFFBB653",
      x"FFFCA62F",
      x"FFFDBE55",
      x"FFFCB344",
      x"FFF79319",
      x"FFF48D15",
      x"FFF18E19",
      x"FFED942A",
      x"FFE9841B",
      x"FFF08814",
      x"FFF29017",
      x"FFF48D16",
      x"FFF39218",
      x"FFE77A0F",
      x"FFDA6F10",
      x"FFD06610",
      x"FFD87117",
      x"FFD87318",
      x"FFDD7E20",
      x"FFDA771B",
      x"FFD67117",
      x"FFD9781C",
      x"FFD0731B",
      x"FFCE721C",
      x"FFC7711E",
      x"FFD37D22",
      x"FFD58225",
      x"FFD57D20",
      x"FFDE8623",
      x"FFE39330",
      x"FFDE9136",
      x"FFD89139",
      x"FFD7913E",
      x"FFD58F3A",
      x"FFD18A38",
      x"FFCE8431",
      x"FFCF8331",
      x"FFDB9244",
      x"FFD88B36",
      x"FFD6852E",
      x"FFD2852B",
      x"FFE68A30",
      x"FFE99138",
      x"FFE5862A",
      x"FFEA9032",
      x"FFEB9438",
      x"FFE99139",
      x"FFEE953F",
      x"FFEF983F",
      x"FFEB943F",
      x"FFF19C45",
      x"FFF4A554",
      x"FFF2A554",
      x"FFEB9A48",
      x"FFE7913F",
      x"FFE58D3D",
      x"FFEEA357",
      x"FFEB9C4B",
      x"FFF0A958",
      x"FFF3AC4C",
      x"FFF9B24E",
      x"FFFAA32C",
      x"FFFDB648",
      x"FFFEBC4E",
      x"FFF89D21",
      x"FFF68F17",
      x"FFF49319",
      x"FFEF982B",
      x"FFEB8B21",
      x"FFF28E19",
      x"FFF08F1A",
      x"FFF38C14",
      x"FFF28B12",
      x"FFE87C0E",
      x"FFDF7513",
      x"FFD1690F",
      x"FFD77218",
      x"FFD57117",
      x"FFD67118",
      x"FFD67118",
      x"FFD67015",
      x"FFD67117",
      x"FFD06F18",
      x"FFD0751D",
      x"FFCD741D",
      x"FFD17921",
      x"FFD58227",
      x"FFD67E21",
      x"FFDD8623",
      x"FFE5912C",
      x"FFDD9233",
      x"FFD68B33",
      x"FFD8923E",
      x"FFD69039",
      x"FFD08936",
      x"FFCF8836",
      x"FFD08736",
      x"FFD88D3D",
      x"FFD98F3E",
      x"FFD68631",
      x"FFD28429",
      x"FFE78C32",
      x"FFE7903A",
      x"FFE5862C",
      x"FFEA8F31",
      x"FFE7882A",
      x"FFEA9039",
      x"FFEC9139",
      x"FFEB8E35",
      x"FFED9744",
      x"FFEC943D",
      x"FFF1A24F",
      x"FFF2A554",
      x"FFEC9C4C",
      x"FFE79241",
      x"FFE58F42",
      x"FFED9B4D",
      x"FFED9D4F",
      x"FFEDA24B",
      x"FFF1AB51",
      x"FFF8B250",
      x"FFFAA62F",
      x"FFFCAD36",
      x"FFFDBD52",
      x"FFFAA72D",
      x"FFF78F15",
      x"FFF79C23",
      x"FFF29A28",
      x"FFED9128",
      x"FFEF8F1E",
      x"FFF49419",
      x"FFF08A14",
      x"FFF49419",
      x"FFE88114",
      x"FFE47F15",
      x"FFD2650D",
      x"FFD26A13",
      x"FFD97518",
      x"FFD56C15",
      x"FFD57217",
      x"FFDB771B",
      x"FFD56E14",
      x"FFD37018",
      x"FFCE711A",
      x"FFD57E23",
      x"FFD47D23",
      x"FFD48226",
      x"FFD88023",
      x"FFDA8220",
      x"FFE38D28",
      x"FFDF9332",
      x"FFD88C34",
      x"FFD68E3A",
      x"FFD6903A",
      x"FFCF8936",
      x"FFD28A37",
      x"FFCE8536",
      x"FFD88E3F",
      x"FFDA903F",
      x"FFD4842E",
      x"FFD1832C",
      x"FFE88E33",
      x"FFE98E36",
      x"FFE4862C",
      x"FFE78B2C",
      x"FFEA8D30",
      x"FFE98B31",
      x"FFEC933B",
      x"FFEB8F36",
      x"FFED9845",
      x"FFEA913A",
      x"FFEF9F4D",
      x"FFF4A95D",
      x"FFED9C4E",
      x"FFE89341",
      x"FFE69247",
      x"FFEA9649",
      x"FFEE9F4F",
      x"FFEB9A40",
      x"FFEEA650",
      x"FFF4AD4E",
      x"FFF8A530",
      x"FFFCA92B",
      x"FFFDB950",
      x"FFFBB042",
      x"FFF98E13",
      x"FFF79F29",
      x"FFF49F2C",
      x"FFEC9228",
      x"FFEB8C21",
      x"FFF28D14",
      x"FFED8310",
      x"FFF18C12",
      x"FFE87C11",
      x"FFE27910",
      x"FFD5690E",
      x"FFD36A12",
      x"FFD87315",
      x"FFD26813",
      x"FFD77218",
      x"FFD87418",
      x"FFD56F16",
      x"FFD5771C",
      x"FFD0731B",
      x"FFD37920",
      x"FFD68024",
      x"FFD47F23",
      x"FFD68024",
      x"FFDB8222",
      x"FFE18C28",
      x"FFE29838",
      x"FFD88D36",
      x"FFD58D3C",
      x"FFD68F3A",
      x"FFD18937",
      x"FFD28A37",
      x"FFCD8434",
      x"FFD68A39",
      x"FFDC9341",
      x"FFD88A34",
      x"FFD18229",
      x"FFE88B30",
      x"FFE5872D",
      x"FFE78B30",
      x"FFE6892D",
      x"FFEC9132",
      x"FFEA8F33",
      x"FFED953A",
      x"FFEC9036",
      x"FFEB923D",
      x"FFE98F3A",
      x"FFF09E4A",
      x"FFF2A85B",
      x"FFF0A051",
      x"FFEB9745",
      x"FFE69346",
      x"FFE89140",
      x"FFEFA051",
      x"FFEEA04A",
      x"FFECA049",
      x"FFF0A647",
      x"FFF6A633",
      x"FFFBAB2F",
      x"FFFCAF3C",
      x"FFFBB54B",
      x"FFF9971E",
      x"FFF8981D",
      x"FFF59F2A",
      x"FFF09627",
      x"FFED8E23",
      x"FFF2941B",
      x"FFED7D0B",
      x"FFED7F0C",
      x"FFE77A0E",
      x"FFE57F12",
      x"FFD76A0C",
      x"FFD16811",
      x"FFD97215",
      x"FFCE6010",
      x"FFD77116",
      x"FFD66E14",
      x"FFD46B11",
      x"FFD4741B",
      x"FFD0711A",
      x"FFCD761E",
      x"FFD47E22",
      x"FFD58023",
      x"FFD78024",
      x"FFD98221",
      x"FFE08928",
      x"FFE39837",
      x"FFD68933",
      x"FFD58D3B",
      x"FFD6913E",
      x"FFD08835",
      x"FFD18937",
      x"FFCF8735",
      x"FFD38836",
      x"FFDA903E",
      x"FFD88D35",
      x"FFD38429",
      x"FFEA8F34",
      x"FFE98A2F",
      x"FFE88E33",
      x"FFE5892E",
      x"FFEB8F30",
      x"FFEB9034",
      x"FFEC9237",
      x"FFEA8F36",
      x"FFE88A31",
      x"FFE98F3B",
      x"FFEE9B46",
      x"FFF2A75B",
      x"FFF0A355",
      x"FFEC9E50",
      x"FFE79040",
      x"FFE48A3A",
      x"FFEB9849",
      x"FFEFA552",
      x"FFEB9B41",
      x"FFEAA047",
      x"FFF4A537",
      x"FFF9AB37",
      x"FFFDB340",
      x"FFFCB64E",
      x"FFFAA12C",
      x"FFF79015",
      x"FFF69C26",
      x"FFF19726",
      x"FFEF9226",
      x"FFF09322",
      x"FFEF8411",
      x"FFEB7A09",
      x"FFE6750B",
      x"FFE78315",
      x"FFD86D10",
      x"FFD16A12",
      x"FFD87215",
      x"FFD0630F",
      x"FFD87213",
      x"FFD46D13",
      x"FFD26B13",
      x"FFD27018",
      x"FFCD6E18",
      x"FFD2791F",
      x"FFD37C24",
      x"FFD47F22",
      x"FFD78226",
      x"FFDB8121",
      x"FFDF8927",
      x"FFE49A37",
      x"FFD98D33",
      x"FFD78F40",
      x"FFD58C38",
      x"FFD38D3B",
      x"FFD08736",
      x"FFCF8634",
      x"FFD28734",
      x"FFDB913F",
      x"FFD98D37",
      x"FFD5862B",
      x"FFE6892E",
      x"FFEA8C2F",
      x"FFE98D31",
      x"FFE4842A",
      x"FFE78A2D",
      x"FFEB8E30",
      x"FFEB8F35",
      x"FFEB8F35",
      x"FFE98C32",
      x"FFEB933F",
      x"FFEA933D",
      x"FFF2A65C",
      x"FFF2A759",
      x"FFED9E4D",
      x"FFE99545",
      x"FFE3893A",
      x"FFE9913F",
      x"FFF0A654",
      x"FFEC9C43",
      x"FFE89943",
      x"FFF09F37",
      x"FFF7A736",
      x"FFFDB543",
      x"FFFBB446",
      x"FFFBAA3A",
      x"FFF89318",
      x"FFF69E25",
      x"FFF29220",
      x"FFF1992A",
      x"FFF39723",
      x"FFEC8512",
      x"FFE9780B",
      x"FFE4750C",
      x"FFE58113",
      x"FFD4620D",
      x"FFCF6812",
      x"FFD87217",
      x"FFCF6511",
      x"FFD86F12",
      x"FFD97417",
      x"FFD26C12",
      x"FFD16F18",
      x"FFCE6F19",
      x"FFD27920",
      x"FFD37C23",
      x"FFD58023",
      x"FFD88324",
      x"FFDA8122",
      x"FFDE8624",
      x"FFE59937",
      x"FFDC933B",
      x"FFD99243",
      x"FFD58D3A",
      x"FFD18837",
      x"FFD1842D",
      x"FFD08835",
      x"FFD08635",
      x"FFDA903E",
      x"FFD98D36",
      x"FFD7882D",
      x"FFEA8A30",
      x"FFEB8C2F",
      x"FFEB9033",
      x"FFE98B2F",
      x"FFE28327",
      x"FFE98B2C",
      x"FFE88C2F",
      x"FFEA8D31",
      x"FFE9892E",
      x"FFE9903A",
      x"FFE88F3A",
      x"FFF2A454",
      x"FFF2A656",
      x"FFF1A04E",
      x"FFEC9C4D",
      x"FFE58E3E",
      x"FFE68D3E",
      x"FFED9D4B",
      x"FFEFA552",
      x"FFEB993E",
      x"FFED9C3A",
      x"FFF5A02D",
      x"FFFCB84C",
      x"FFFBB13D",
      x"FFFCB144",
      x"FFF9951A",
      x"FFF89F21",
      x"FFF2921E",
      x"FFF29928",
      x"FFF29721",
      x"FFED8913",
      x"FFE97E0F",
      x"FFE77A0F",
      x"FFE17B13",
      x"FFD3600A",
      x"FFCE6510",
      x"FFD67116",
      x"FFD06813",
      x"FFD77013",
      x"FFD77115",
      x"FFD26D13",
      x"FFCE6B16",
      x"FFCD6E18",
      x"FFD2761E",
      x"FFD17921",
      x"FFD67F22",
      x"FFD68124",
      x"FFDC8626",
      x"FFDE8523",
      x"FFE49533",
      x"FFDA8D33",
      x"FFD89244",
      x"FFD58C3A",
      x"FFD18938",
      x"FFD08530",
      x"FFCE8634",
      x"FFD18635",
      x"FFD98E3A",
      x"FFDC913B",
      x"FFD6892E",
      x"FFEA8E2F",
      x"FFE98D30",
      x"FFEB8E30",
      x"FFE98B2E",
      x"FFE48425",
      x"FFEC9131",
      x"FFEB8C2D",
      x"FFEC9133",
      x"FFEA8E33",
      x"FFEC933A",
      x"FFE9913B",
      x"FFF1A451",
      x"FFF3A857",
      x"FFF1A454",
      x"FFED9B47",
      x"FFE5903E",
      x"FFE38738",
      x"FFEB9947",
      x"FFF2AA56",
      x"FFEB9537",
      x"FFE9983D",
      x"FFF2A032",
      x"FFFCB547",
      x"FFFCAF3A",
      x"FFFBAE3D",
      x"FFFBA125",
      x"FFF69C22",
      x"FFF29320",
      x"FFF08E1B",
      x"FFF09526",
      x"FFEC8614",
      x"FFE5790C",
      x"FFE4770F",
      x"FFE37E15",
      x"FFD6660D",
      x"FFD06611",
      x"FFD66F15",
      x"FFCF6511",
      x"FFD66E12",
      x"FFD56C12",
      x"FFD36C13",
      x"FFCD6813",
      x"FFD06F19",
      x"FFD2771F",
      x"FFD37921",
      x"FFD47B20",
      x"FFD68022",
      x"FFDA8122",
      x"FFDF8522",
      x"FFE59733",
      x"FFDC8F32",
      x"FFD78E3D",
      x"FFD68D3B",
      x"FFD18A38",
      x"FFCD812F",
      x"FFCF8530",
      x"FFCF8431",
      x"FFDB8E39",
      x"FFDC913C",
      x"FFD88C32",
      x"FFEA8D33",
      x"FFE98E30",
      x"FFE88B2E",
      x"FFE89036",
      x"FFE38328",
      x"FFEA8C2B",
      x"FFEB8F31",
      x"FFE98C30",
      x"FFEA8C2F",
      x"FFEB9135",
      x"FFE78C36",
      x"FFEF9C44",
      x"FFF3A756",
      x"FFF2A553",
      x"FFEE9A43",
      x"FFE99644",
      x"FFE48C3C",
      x"FFEA9240",
      x"FFEFA453",
      x"FFEA9337",
      x"FFE89438",
      x"FFED9832",
      x"FFF5A93B",
      x"FFFCB446",
      x"FFFBAC32",
      x"FFFCA92E",
      x"FFFAA628",
      x"FFF59B27",
      x"FFF39421",
      x"FFF19B2B",
      x"FFE97F10",
      x"FFE5760B",
      x"FFE1710B",
      x"FFE57F15",
      x"FFD5660D",
      x"FFD16912",
      x"FFD76F14",
      x"FFCE6410",
      x"FFD46D10",
      x"FFD77015",
      x"FFD36D14",
      x"FFCC6712",
      x"FFD06F18",
      x"FFD1751D",
      x"FFD37A21",
      x"FFD37C22",
      x"FFD68123",
      x"FFDB8422",
      x"FFE18825",
      x"FFE69A36",
      x"FFDB8C30",
      x"FFD68D3B",
      x"FFD68D3B",
      x"FFD28A3A",
      x"FFCB802C",
      x"FFCE8330",
      x"FFD28837",
      x"FFD98B37",
      x"FFDD943F",
      x"FFD6872B",
      x"FFEA8F31",
      x"FFE98A2E",
      x"FFE98C30",
      x"FFEA8F34",
      x"FFE68A30",
      x"FFE78729",
      x"FFEA8D2C",
      x"FFEA8B2F",
      x"FFEA8C30",
      x"FFE88A2F",
      x"FFEA9037",
      x"FFED953D",
      x"FFF3A853",
      x"FFF3A85A",
      x"FFF09F4C",
      x"FFEC9944",
      x"FFE58E3F",
      x"FFE8903F",
      x"FFEB9A47",
      x"FFEC9A41",
      x"FFE78D33",
      x"FFEA9637",
      x"FFF3A131",
      x"FFFCB647",
      x"FFFCAD39",
      x"FFFBA52C",
      x"FFFBA221",
      x"FFF4941E",
      x"FFF39520",
      x"FFF19B2D",
      x"FFE88113",
      x"FFE57309",
      x"FFE06B08",
      x"FFE47E15",
      x"FFD86B0F",
      x"FFD36A14",
      x"FFD56A13",
      x"FFCD6310",
      x"FFD3690E",
      x"FFD46C12",
      x"FFD57116",
      x"FFC9610F",
      x"FFCF6C15",
      x"FFD4761C",
      x"FFD67C22",
      x"FFD47B20",
      x"FFD98023",
      x"FFDB8223",
      x"FFE18A26",
      x"FFE99C3A",
      x"FFDD9032",
      x"FFD58B38",
      x"FFD48B3A",
      x"FFD38B3C",
      x"FFCD8332",
      x"FFCC8432",
      x"FFD18634",
      x"FFD88A35",
      x"FFDF953F",
      x"FFDA8C2F",
      x"FFED9435",
      x"FFE58529",
      x"FFE4872F",
      x"FFE88C30",
      x"FFE78A2C",
      x"FFE48124",
      x"FFEC9231",
      x"FFEA8D2F",
      x"FFED9134",
      x"FFE8882B",
      x"FFEC933B",
      x"FFED963E",
      x"FFF2A34E",
      x"FFF3AA5B",
      x"FFF1A04F",
      x"FFEC9840",
      x"FFE58C39",
      x"FFE89345",
      x"FFE89242",
      x"FFEC9C47",
      x"FFE78E33",
      x"FFEA9739",
      x"FFEE982B",
      x"FFFBB33F",
      x"FFFBB23F",
      x"FFF9A028",
      x"FFFAA223",
      x"FFF3931D",
      x"FFF59118",
      x"FFF09526",
      x"FFEA8416",
      x"FFE5780C",
      x"FFE16F09",
      x"FFDD7211",
      x"FFD5670D",
      x"FFD46F14",
      x"FFD56A11",
      x"FFD06812",
      x"FFCF620B",
      x"FFD16B10",
      x"FFD67417",
      x"FFC8610F",
      x"FFCE6E17",
      x"FFD57A1F",
      x"FFD87D20",
      x"FFD77E22",
      x"FFD67E20",
      x"FFDC8424",
      x"FFDF8523",
      x"FFE89D38",
      x"FFDF9237",
      x"FFD78E3D",
      x"FFD38A39",
      x"FFD38B3E",
      x"FFD08735",
      x"FFCD8331",
      x"FFCE8433",
      x"FFD78A36",
      x"FFDD923C",
      x"FFDC9036",
      x"FFED9535",
      x"FFEA8E30",
      x"FFE98E30",
      x"FFE6892D",
      x"FFE88D30",
      x"FFE68527",
      x"FFEA8D2D",
      x"FFE98C31",
      x"FFEB8C2D",
      x"FFEC8E2D",
      x"FFEB9037",
      x"FFE88E38",
      x"FFF1A14E",
      x"FFF2A958",
      x"FFF2A453",
      x"FFEC973E",
      x"FFE8903A",
      x"FFE68B38",
      x"FFE78E3D",
      x"FFE68F3A",
      x"FFE89038",
      x"FFE78D30",
      x"FFEB9730",
      x"FFF8A72D",
      x"FFFBAE3C",
      x"FFF8A12A",
      x"FFFAA325",
      x"FFF4931D",
      x"FFF6951B",
      x"FFF39926",
      x"FFEC8B1B",
      x"FFE77E11",
      x"FFE0700C",
      x"FFDB690D",
      x"FFD6670D",
      x"FFD47118",
      x"FFD76E14",
      x"FFD26F14",
      x"FFCC5F0B",
      x"FFD06B12",
      x"FFD36E12",
      x"FFCA630E",
      x"FFCC6A14",
      x"FFD5761B",
      x"FFDC8425",
      x"FFD98224",
      x"FFD78123",
      x"FFDC8525",
      x"FFDF8725",
      x"FFE79A36",
      x"FFDE9236",
      x"FFD48B38",
      x"FFD58B3B",
      x"FFD28633",
      x"FFCE8431",
      x"FFCF8431",
      x"FFD18634",
      x"FFD98B36",
      x"FFDD933E",
      x"FFDE943B",
      x"FFED9230",
      x"FFEB8E31",
      x"FFEA8D30",
      x"FFEA8C2E",
      x"FFE98D2E",
      x"FFE78C30",
      x"FFE7892A",
      x"FFEA8E31",
      x"FFEA8D2F",
      x"FFEA8D2E",
      x"FFEB8E33",
      x"FFEB933B",
      x"FFED993F",
      x"FFF2A651",
      x"FFF1A351",
      x"FFEF9940",
      x"FFEA9139",
      x"FFE48834",
      x"FFEA9241",
      x"FFE78E3B",
      x"FFE99640",
      x"FFE68B30",
      x"FFEA9431",
      x"FFF3A12F",
      x"FFFAAE3A",
      x"FFFAA834",
      x"FFFAA627",
      x"FFF69920",
      x"FFF3931C",
      x"FFF5A02E",
      x"FFEF901D",
      x"FFEA8314",
      x"FFE47A10",
      x"FFD8650A",
      x"FFD6690D",
      x"FFD47017",
      x"FFD66D14",
      x"FFD06C14",
      x"FFC85B0B",
      x"FFD47113",
      x"FFCE660F",
      x"FFC65F0E",
      x"FFCC6812",
      x"FFD6771D",
      x"FFE08928",
      x"FFDD8724",
      x"FFD98425",
      x"FFDE8926",
      x"FFDF8724",
      x"FFE79937",
      x"FFDE9034",
      x"FFD28732",
      x"FFD18332",
      x"FFD48734",
      x"FFD28837",
      x"FFD38735",
      x"FFD1822F",
      x"FFD98B35",
      x"FFE09740",
      x"FFDE963C",
      x"FFE68828",
      x"FFEB8C2D",
      x"FFEA8D2C",
      x"FFEA8F30",
      x"FFE7882B",
      x"FFE9892A",
      x"FFE7892B",
      x"FFE78729",
      x"FFE98C2F",
      x"FFEC9034",
      x"FFE78528",
      x"FFEC933A",
      x"FFEB933B",
      x"FFF1A350",
      x"FFF0A251",
      x"FFF19E48",
      x"FFEC953F",
      x"FFE48936",
      x"FFE7903E",
      x"FFE68C3A",
      x"FFE8933C",
      x"FFE79039",
      x"FFE68E2D",
      x"FFF09F34",
      x"FFF7A834",
      x"FFFAAB34",
      x"FFFAA82E",
      x"FFF89F23",
      x"FFF1911E",
      x"FFF5A02C",
      x"FFF0921D",
      x"FFE98515",
      x"FFE67F11",
      x"FFDC6F0F",
      x"FFD7670D",
      x"FFD57017",
      x"FFD46A13",
      x"FFD36E13",
      x"FFC9590A",
      x"FFD56F12",
      x"FFD06A11",
      x"FFCA620D",
      x"FFCD6A13",
      x"FFD77A1D",
      x"FFDF8825",
      x"FFE08C28",
      x"FFDB8624",
      x"FFDD8927",
      x"FFE38E2A",
      x"FFE79C39",
      x"FFDD8D2E",
      x"FFD78E3D",
      x"FFD48836",
      x"FFD88C38",
      x"FFD18735",
      x"FFD48836",
      x"FFD48632",
      x"FFD88A34",
      x"FFE09641",
      x"FFDD923B",
      x"FFEC8E2D",
      x"FFEB8C2C",
      x"FFE9882A",
      x"FFEA8D2E",
      x"FFE8892B",
      x"FFE88C2D",
      x"FFE58728",
      x"FFE98D2D",
      x"FFE68729",
      x"FFEC8E31",
      x"FFE98A2C",
      x"FFE98F36",
      x"FFEA923D",
      x"FFF1A24C",
      x"FFF0A04F",
      x"FFF09D48",
      x"FFE9933C",
      x"FFE58B35",
      x"FFE68E3C",
      x"FFE88E3A",
      x"FFE5862E",
      x"FFE68B32",
      x"FFE5892B",
      x"FFED982D",
      x"FFF4A432",
      x"FFF8A82E",
      x"FFF7A429",
      x"FFF8A226",
      x"FFEF8F20",
      x"FFF49D2C",
      x"FFF29822",
      x"FFEB8917",
      x"FFE68012",
      x"FFDD6C0C",
      x"FFD66109",
      x"FFD46E14",
      x"FFCD5E0D",
      x"FFD26A11",
      x"FFCA5E0B",
      x"FFD36B0F",
      x"FFD36C11",
      x"FFCC660E",
      x"FFCD6A13",
      x"FFD4761A",
      x"FFE18D2A",
      x"FFDF8C29",
      x"FFDC8C28",
      x"FFDD8A28",
      x"FFE28D2A",
      x"FFE89C39",
      x"FFE09436",
      x"FFD9903B",
      x"FFD28939",
      x"FFD78A39",
      x"FFD38835",
      x"FFD28532",
      x"FFD68934",
      x"FFDB8D36",
      x"FFDE943E",
      x"FFDB933B",
      x"FFED902F",
      x"FFEC902F",
      x"FFEA8C2F",
      x"FFEC9131",
      x"FFE78425",
      x"FFE98D2E",
      x"FFE48325",
      x"FFE58729",
      x"FFEA8E2F",
      x"FFEC9133",
      x"FFEA8F31",
      x"FFEB9034",
      x"FFE99139",
      x"FFF19D44",
      x"FFF1A04C",
      x"FFF09F4A",
      x"FFEC933C",
      x"FFE8903B",
      x"FFE78D38",
      x"FFE88F3D",
      x"FFE78A32",
      x"FFE38329",
      x"FFE48528",
      x"FFE8902C",
      x"FFF1A438",
      x"FFF6A52C",
      x"FFF8A324",
      x"FFFAA729",
      x"FFEF9323",
      x"FFF39D2A",
      x"FFF49D26",
      x"FFEE8F1A",
      x"FFE98213",
      x"FFE07510",
      x"FFD66309",
      x"FFD67114",
      x"FFCD5C0D",
      x"FFD16810",
      x"FFC85B0C",
      x"FFD16A0F",
      x"FFCD670E",
      x"FFC7620E",
      x"FFCD6A11",
      x"FFD6771A",
      x"FFE08B28",
      x"FFE1902D",
      x"FFDD8B27",
      x"FFDC8927",
      x"FFE18C28",
      x"FFE49634",
      x"FFE2963B",
      x"FFD58B34",
      x"FFD58C39",
      x"FFD58A3B",
      x"FFD38532",
      x"FFD28534",
      x"FFDC8F3E",
      x"FFDF933D",
      x"FFDC8C36",
      x"FFDA923E",
      x"FFED8F2B",
      x"FFEB8B2B",
      x"FFE88629",
      x"FFEA8E2F",
      x"FFE68425",
      x"FFE78727",
      x"FFE78828",
      x"FFE18023",
      x"FFE8892A",
      x"FFE98E30",
      x"FFEA8C2C",
      x"FFEA8B2D",
      x"FFE88D34",
      x"FFEC963B",
      x"FFF19E4A",
      x"FFEF9E48",
      x"FFED953A",
      x"FFEA953F",
      x"FFE68B33",
      x"FFE88D3A",
      x"FFE78A31",
      x"FFE58930",
      x"FFE4842A",
      x"FFE48424",
      x"FFED9B33",
      x"FFF3A230",
      x"FFF6A223",
      x"FFFAA729",
      x"FFF09726",
      x"FFF19A28",
      x"FFF59C22",
      x"FFF1951F",
      x"FFEA8111",
      x"FFE0750F",
      x"FFD9690C",
      x"FFD77316",
      x"FFCF6210",
      x"FFD26C14",
      x"FFC9590B",
      x"FFD26A0E",
      x"FFCE680F",
      x"FFCB6911",
      x"FFCE6B11",
      x"FFD97C1D",
      x"FFE38F2B",
      x"FFE0912E",
      x"FFDC8A27",
      x"FFDA8A29",
      x"FFE2902A",
      x"FFE39633",
      x"FFDF9336",
      x"FFD88C39",
      x"FFD58A38",
      x"FFD58937",
      x"FFD68935",
      x"FFD28434",
      x"FFD88A37",
      x"FFDD8F3A",
      x"FFE1943E",
      x"FFDA8F3C",
      x"FFED902B",
      x"FFEB8926",
      x"FFE88527",
      x"FFE98929",
      x"FFE58427",
      x"FFE58124",
      x"FFE38224",
      x"FFE17F23",
      x"FFE88A2A",
      x"FFE88A2D",
      x"FFE88626",
      x"FFE78326",
      x"FFE88C33",
      x"FFE88F35",
      x"FFF09D46",
      x"FFEF9E49",
      x"FFED953E",
      x"FFEA933C",
      x"FFE68930",
      x"FFE88D3A",
      x"FFE78B35",
      x"FFE1842C",
      x"FFE4882E",
      x"FFE37F21",
      x"FFE9922B",
      x"FFF1A034",
      x"FFF49F21",
      x"FFF9A92D",
      x"FFF29823",
      x"FFEB8E20",
      x"FFF3951B",
      x"FFF2951C",
      x"FFEA800F",
      x"FFE17911",
      x"FFDE7815",
      x"FFD66F13",
      x"FFCD6211",
      x"FFD46E14",
      x"FFC85B0B",
      x"FFD26D10",
      x"FFCF680F",
      x"FFCD6910",
      x"FFCD6A12",
      x"FFDB7F1D",
      x"FFE28F2B",
      x"FFE09330",
      x"FFDE8E2B",
      x"FFDA8728",
      x"FFE39530",
      x"FFE2912F",
      x"FFDF9338",
      x"FFD98E38",
      x"FFD68A37",
      x"FFD78939",
      x"FFD88B38",
      x"FFD48834",
      x"FFD98C36",
      x"FFDD923C",
      x"FFDF923E",
      x"FFDB8F3B",
      x"FFEC8822",
      x"FFEB8A26",
      x"FFE98827",
      x"FFE98828",
      x"FFE68527",
      x"FFE58425",
      x"FFE78829",
      x"FFE27E21",
      x"FFE78628",
      x"FFE88C2B",
      x"FFEC8F2E",
      x"FFEA8627",
      x"FFE7892D",
      x"FFE78B31",
      x"FFEF993F",
      x"FFEF9B45",
      x"FFED9236",
      x"FFEA9035",
      x"FFE58A32",
      x"FFE68835",
      x"FFE78934",
      x"FFE2812A",
      x"FFDF812A",
      x"FFE0781E",
      x"FFE58A27",
      x"FFEE9A33",
      x"FFF3A027",
      x"FFF8AB32",
      x"FFF39B27",
      x"FFEB8B1D",
      x"FFEE8B15",
      x"FFF18D13",
      x"FFED8814",
      x"FFE1760E",
      x"FFDB7614",
      x"FFD67016",
      x"FFCE6413",
      x"FFD67316",
      x"FFC7580A",
      x"FFD16A0F",
      x"FFCE660D",
      x"FFCC6A10",
      x"FFCB6910",
      x"FFDC821F",
      x"FFE2902C",
      x"FFDF8F2D",
      x"FFDB8F2E",
      x"FFDA8A2A",
      x"FFE2932F",
      x"FFE28F2D",
      x"FFE09437",
      x"FFD88C37",
      x"FFD58A38",
      x"FFD88A3A",
      x"FFD98E3B",
      x"FFD78936",
      x"FFDB8D37",
      x"FFDD903C",
      x"FFDC8F3A",
      x"FFDA852A",
      x"FFE7811D",
      x"FFEB8925",
      x"FFEA8926",
      x"FFE78629",
      x"FFE98829",
      x"FFE68022",
      x"FFE98828",
      x"FFE88A2A",
      x"FFE48020",
      x"FFE88A2C",
      x"FFED9231",
      x"FFEB8B29",
      x"FFE78B30",
      x"FFE5862E",
      x"FFEE963B",
      x"FFF19D45",
      x"FFEE963C",
      x"FFEB8C2F",
      x"FFE78D37",
      x"FFE58834",
      x"FFE68A35",
      x"FFE68B35",
      x"FFDD7C27",
      x"FFE17A1F",
      x"FFE08020",
      x"FFEA932E",
      x"FFF19E2C",
      x"FFF6A82F",
      x"FFF49D2A",
      x"FFEC8B1C",
      x"FFEA8313",
      x"FFF39016",
      x"FFEE8F19",
      x"FFE1760F",
      x"FFDC6E0F",
      x"FFD36B10",
      x"FFD06614",
      x"FFD77116",
      x"FFC8590B",
      x"FFD0680D",
      x"FFCF680E",
      x"FFCD6A10",
      x"FFC8640E",
      x"FFDB811F",
      x"FFE28E29",
      x"FFE0922F",
      x"FFDB9030",
      x"FFD88C2C",
      x"FFDF9230",
      x"FFE3922F",
      x"FFDF9133",
      x"FFD88C38",
      x"FFD58B3A",
      x"FFDB8F3F",
      x"FFDB8E3B",
      x"FFD98B34",
      x"FFD98A34",
      x"FFDF9642",
      x"FFDC903B",
      x"FFDD8729",
      x"FFE9821C",
      x"FFEE9127",
      x"FFED8A27",
      x"FFEA8B2C",
      x"FFE98627",
      x"FFEA882A",
      x"FFE98627",
      x"FFE98B2A",
      x"FFE88928",
      x"FFE98726",
      x"FFEB8F2E",
      x"FFEF9331",
      x"FFEC8F31",
      x"FFEB8D32",
      x"FFEC8D31",
      x"FFEF9B42",
      x"FFED963B",
      x"FFEB8E30",
      x"FFE9913A",
      x"FFE58830",
      x"FFE78D3A",
      x"FFE68932",
      x"FFE0802C",
      x"FFE37F23",
      x"FFDC7217",
      x"FFE58A27",
      x"FFEF9A2D",
      x"FFF4A327",
      x"FFF7A631",
      x"FFED8D1D",
      x"FFE87E11",
      x"FFF29017",
      x"FFF09119",
      x"FFE57C10",
      x"FFDA6F0E",
      x"FFD36A13",
      x"FFD06513",
      x"FFD87418",
      x"FFC95E0E",
      x"FFD56F0F",
      x"FFCB640D",
      x"FFCE6C12",
      x"FFCB660E",
      x"FFD97E1D",
      x"FFE2912C",
      x"FFE09633",
      x"FFDA8E31",
      x"FFD6892C",
      x"FFDD8E2D",
      x"FFE39333",
      x"FFDE9133",
      x"FFDA903D",
      x"FFD3893B",
      x"FFD98D3B",
      x"FFDB8D39",
      x"FFDA8A31",
      x"FFD98A34",
      x"FFDE943D",
      x"FFDE9644",
      x"FFDF8E36",
      x"FFEA861F",
      x"FFEE9029",
      x"FFEF932D",
      x"FFEA8927",
      x"FFE68224",
      x"FFE98B2B",
      x"FFE9892A",
      x"FFE7892B",
      x"FFE68324",
      x"FFE88825",
      x"FFE88A2C",
      x"FFED8F2F",
      x"FFEC9234",
      x"FFEB9134",
      x"FFEB9031",
      x"FFF1A04A",
      x"FFEE9941",
      x"FFEB9035",
      x"FFEA913A",
      x"FFE48731",
      x"FFE58531",
      x"FFE78933",
      x"FFE3822C",
      x"FFE17C21",
      x"FFDE7118",
      x"FFE07F20",
      x"FFEB942D",
      x"FFF29D22",
      x"FFF6A832",
      x"FFF0901D",
      x"FFE67C12",
      x"FFED8A17",
      x"FFEF911B",
      x"FFE67E0F",
      x"FFDB7514",
      x"FFD0610D",
      x"FFCD6212",
      x"FFD87619",
      x"FFCC600F",
      x"FFD56F12",
      x"FFCD670E",
      x"FFCD6B11",
      x"FFCC660F",
      x"FFDA7E1D",
      x"FFE39430",
      x"FFE09636",
      x"FFD88C2F",
      x"FFD4872B",
      x"FFDB8C2B",
      x"FFE08E2C",
      x"FFDF9031",
      x"FFD98C36",
      x"FFD58B39",
      x"FFDB8C3B",
      x"FFDB8D3B",
      x"FFDD9039",
      x"FFDD903C",
      x"FFDF943E",
      x"FFDC9541",
      x"FFDD8C36",
      x"FFEB8821",
      x"FFEC8C24",
      x"FFEE8D28",
      x"FFEC8E2B",
      x"FFEB8929",
      x"FFE98728",
      x"FFE7882A",
      x"FFE88A2C",
      x"FFE58324",
      x"FFE78624",
      x"FFE58627",
      x"FFED8F2D",
      x"FFEC8F2E",
      x"FFED9539",
      x"FFEC9134",
      x"FFF3A34D",
      x"FFED983F",
      x"FFEA9136",
      x"FFEA923A",
      x"FFE68B36",
      x"FFE78B35",
      x"FFE78A33",
      x"FFE4852E",
      x"FFE5862C",
      x"FFDF7219",
      x"FFE17F22",
      x"FFEA9330",
      x"FFF19B24",
      x"FFF5A42D",
      x"FFF39720",
      x"FFEB8717",
      x"FFE88217",
      x"FFEF8F1B",
      x"FFE78010",
      x"FFDB7313",
      x"FFD36610",
      x"FFCC5D0F",
      x"FFD87219",
      x"FFCE610F",
      x"FFD2690F",
      x"FFCD670F",
      x"FFCD6810",
      x"FFCA660E",
      x"FFDA801F",
      x"FFDE8D2A",
      x"FFD99030",
      x"FFD58B2E",
      x"FFD2832A",
      x"FFD78729",
      x"FFDF8E2E",
      x"FFE19438",
      x"FFD88A34",
      x"FFD78C3B",
      x"FFD98D3A",
      x"FFDA8B36",
      x"FFDC8E37",
      x"FFDD8F36",
      x"FFDE953D",
      x"FFDC923D",
      x"FFDA862F",
      x"FFED8E26",
      x"FFEF8F26",
      x"FFEF8E26",
      x"FFEC8D2B",
      x"FFEC8D29",
      x"FFE88424",
      x"FFE68427",
      x"FFE58428",
      x"FFE58525",
      x"FFE48121",
      x"FFE6872B",
      x"FFEB8D2C",
      x"FFEC8D2C",
      x"FFEC9336",
      x"FFEA8F34",
      x"FFF2A149",
      x"FFED9845",
      x"FFEB943A",
      x"FFE9913D",
      x"FFE58B36",
      x"FFE78B37",
      x"FFE98E37",
      x"FFE68732",
      x"FFE68B31",
      x"FFE37920",
      x"FFE07B22",
      x"FFE78C28",
      x"FFED9422",
      x"FFF49F25",
      x"FFF39924",
      x"FFE98416",
      x"FFE67D14",
      x"FFED901D",
      x"FFE78516",
      x"FFDB7616",
      x"FFCF620F",
      x"FFCE5F0F",
      x"FFD57019",
      x"FFCF650F",
      x"FFD2690E",
      x"FFD06B10",
      x"FFCF6E12",
      x"FFD06A0F",
      x"FFDB7F1C",
      x"FFE08D28",
      x"FFDC9232",
      x"FFD68B30",
      x"FFD2842B",
      x"FFD7892D",
      x"FFD9892A",
      x"FFE19438",
      x"FFD88835",
      x"FFD68B3B",
      x"FFDB8E3C",
      x"FFDB8E37",
      x"FFDB8C35",
      x"FFE0953C",
      x"FFDF9842",
      x"FFDD9341",
      x"FFDB872F",
      x"FFEA8820",
      x"FFED8E28",
      x"FFEE8F28",
      x"FFEA8B28",
      x"FFED8E2A",
      x"FFE98523",
      x"FFE98928",
      x"FFE58122",
      x"FFE48225",
      x"FFE38121",
      x"FFE5872A",
      x"FFE98A2A",
      x"FFED8E2C",
      x"FFEE9638",
      x"FFEB8E33",
      x"FFF1A049",
      x"FFED9840",
      x"FFED9943",
      x"FFEC9944",
      x"FFE38931",
      x"FFE88D38",
      x"FFE88C33",
      x"FFE78B33",
      x"FFE5882F",
      x"FFE17A21",
      x"FFDF761D",
      x"FFE68C2B",
      x"FFEC9322",
      x"FFF39920",
      x"FFF09320",
      x"FFED9120",
      x"FFE67B10",
      x"FFEC8D1E",
      x"FFE88817",
      x"FFDC7614",
      x"FFCF5F0E",
      x"FFD05F0F",
      x"FFD56E19",
      x"FFCF6612",
      x"FFD2670E",
      x"FFD26F12",
      x"FFD16D10",
      x"FFCE670E",
      x"FFDD831E",
      x"FFE18E2A",
      x"FFDC9232",
      x"FFD4892E",
      x"FFD2852C",
      x"FFD7852A",
      x"FFD88427",
      x"FFDE9032",
      x"FFD88834",
      x"FFD68836",
      x"FFDD9040",
      x"FFDD8C34",
      x"FFDD8E37",
      x"FFDE8F33",
      x"FFE1983F",
      x"FFDC933F",
      x"FFDB8830",
      x"FFE88621",
      x"FFE68120",
      x"FFEA8925",
      x"FFEB8F2D",
      x"FFEA8B2A",
      x"FFEA8927",
      x"FFE88728",
      x"FFE88A2C",
      x"FFE68627",
      x"FFE27E20",
      x"FFE6862A",
      x"FFEB8D2C",
      x"FFEA8C2B",
      x"FFEB9031",
      x"FFE7882D",
      x"FFF09D45",
      x"FFEE9D4A",
      x"FFEC9642",
      x"FFEA9643",
      x"FFE58C38",
      x"FFE88F3D",
      x"FFEA8F39",
      x"FFEB933E",
      x"FFE3872F",
      x"FFE17A20",
      x"FFE0721A",
      x"FFE48829",
      x"FFEC9424",
      x"FFF39C24",
      x"FFEF901E",
      x"FFEF9220",
      x"FFE67D12",
      x"FFE8831A",
      x"FFE98A1B",
      x"FFE07D19",
      x"FFD06410",
      x"FFD57219",
      x"FFD46B16",
      x"FFD26D16",
      x"FFD36B11",
      x"FFD26F12",
      x"FFD27215",
      x"FFCF6A0F",
      x"FFDE8420",
      x"FFE0912A",
      x"FFDC9231",
      x"FFD1842C",
      x"FFD4842A",
      x"FFD8882C",
      x"FFD68227",
      x"FFDE9035",
      x"FFD88935",
      x"FFD78A3B",
      x"FFDD9140",
      x"FFE08F37",
      x"FFDE9236",
      x"FFE09333",
      x"FFE09439",
      x"FFDB903B",
      x"FFD9862D",
      x"FFEC8C22",
      x"FFE47C1B",
      x"FFEC8C29",
      x"FFE9892A",
      x"FFEB8D2D",
      x"FFEA8927",
      x"FFEA8C2C",
      x"FFE68829",
      x"FFE58727",
      x"FFE37F20",
      x"FFE7882A",
      x"FFEA8B29",
      x"FFEC902E",
      x"FFED9233",
      x"FFE98B2E",
      x"FFEE9941",
      x"FFED9C4B",
      x"FFEC9843",
      x"FFE9923B",
      x"FFE1832C",
      x"FFE89242",
      x"FFE88D39",
      x"FFEB9746",
      x"FFE4882F",
      x"FFE0791F",
      x"FFE0761C",
      x"FFE38727",
      x"FFEC9223",
      x"FFF39F27",
      x"FFED8919",
      x"FFEF9826",
      x"FFE78017",
      x"FFE7831C",
      x"FFEA8C1E",
      x"FFE07C18",
      x"FFD26712",
      x"FFD8771C",
      x"FFD26B17",
      x"FFD47019",
      x"FFD1690F",
      x"FFD16C0F",
      x"FFD06E11",
      x"FFD16D0F",
      x"FFDE841D",
      x"FFE3942D",
      x"FFDB9234",
      x"FFD2862C",
      x"FFD5832A",
      x"FFD9882B",
      x"FFD57F25",
      x"FFDD8F37",
      x"FFD78531",
      x"FFD98937",
      x"FFDD8F3C",
      x"FFE09138",
      x"FFE09135",
      x"FFDF9032",
      x"FFDD9035",
      x"FFDA8F3A",
      x"FFDA872D",
      x"FFEB8E26",
      x"FFE98420",
      x"FFEC8C28",
      x"FFEA8C2B",
      x"FFE9892A",
      x"FFEC8E2C",
      x"FFEC8B29",
      x"FFE68526",
      x"FFE68628",
      x"FFE27D1F",
      x"FFE88A2B",
      x"FFEA8D2D",
      x"FFEC8F2D",
      x"FFF09634",
      x"FFEA8C30",
      x"FFEE9A45",
      x"FFEC9947",
      x"FFEE9946",
      x"FFE99641",
      x"FFE48936",
      x"FFE79243",
      x"FFEA9140",
      x"FFE8903F",
      x"FFE58935",
      x"FFDE781F",
      x"FFE0761E",
      x"FFE28326",
      x"FFEB9123",
      x"FFF2A029",
      x"FFEF901E",
      x"FFF19B28",
      x"FFE88519",
      x"FFE17B18",
      x"FFE98B1F",
      x"FFE07E1B",
      x"FFD26610",
      x"FFD7771D",
      x"FFD06919",
      x"FFD47019",
      x"FFD0660F",
      x"FFD16D10",
      x"FFD06F12",
      x"FFD06A0D",
      x"FFE0861F",
      x"FFE1922D",
      x"FFD99133",
      x"FFD38B33",
      x"FFD7872E",
      x"FFD98428",
      x"FFD68124",
      x"FFDA8A2F",
      x"FFD78632",
      x"FFD98938",
      x"FFDD8D39",
      x"FFE0923A",
      x"FFE09337",
      x"FFDF9233",
      x"FFDD9237",
      x"FFDB8F39",
      x"FFDC882E",
      x"FFE78722",
      x"FFE67E1C",
      x"FFEB8926",
      x"FFEB8C2C",
      x"FFE88829",
      x"FFEB8C2B",
      x"FFEB8B29",
      x"FFE88628",
      x"FFE7892A",
      x"FFE0791C",
      x"FFE78929",
      x"FFE8892B",
      x"FFEA8B2B",
      x"FFED9435",
      x"FFEA8E32",
      x"FFEE9843",
      x"FFEE9C4A",
      x"FFEA9541",
      x"FFE8933F",
      x"FFE48B39",
      x"FFE8903F",
      x"FFE8903E",
      x"FFE8903D",
      x"FFE58B37",
      x"FFE07A20",
      x"FFE1761D",
      x"FFDF7D23",
      x"FFE88D21",
      x"FFF2A42D",
      x"FFEF9421",
      x"FFF3A32F",
      x"FFEA891D",
      x"FFE67F18",
      x"FFE7871D",
      x"FFE3811D",
      x"FFD1640E",
      x"FFD6761C",
      x"FFD46A17",
      x"FFD6721A",
      x"FFCF6710",
      x"FFD16E11",
      x"FFD17013",
      x"FFCE690F",
      x"FFDE821C",
      x"FFE2912A",
      x"FFD68A2A",
      x"FFD3872E",
      x"FFD68229",
      x"FFDB882B",
      x"FFD57E25",
      x"FFDA872C",
      x"FFD78631",
      x"FFDA8B3A",
      x"FFDC8B39",
      x"FFDF9038",
      x"FFDF9035",
      x"FFE09537",
      x"FFDF9335",
      x"FFDA8D38",
      x"FFDC892D",
      x"FFE68725",
      x"FFE5801F",
      x"FFE98321",
      x"FFEB8D29",
      x"FFEA8B2B",
      x"FFE98827",
      x"FFEC8E2A",
      x"FFE78729",
      x"FFE7892A",
      x"FFE48022",
      x"FFE68929",
      x"FFE98A2B",
      x"FFEA8D2F",
      x"FFEC9437",
      x"FFE7892D",
      x"FFEE9841",
      x"FFEE9B47",
      x"FFE99543",
      x"FFE89443",
      x"FFE58B38",
      x"FFE99040",
      x"FFEB9547",
      x"FFE88E3B",
      x"FFE68C37",
      x"FFDD751D",
      x"FFE0761C",
      x"FFDD751D",
      x"FFE4831B",
      x"FFEE9B27",
      x"FFEB8F22",
      x"FFF29F2B",
      x"FFEE9022",
      x"FFE58019",
      x"FFE68219",
      x"FFE2821D",
      x"FFD66C14",
      x"FFD6781E",
      x"FFD36A18",
      x"FFD6731A",
      x"FFD16811",
      x"FFD47214",
      x"FFD16D12",
      x"FFCF6A0F",
      x"FFDF851F",
      x"FFE19430",
      x"FFD89033",
      x"FFD4872D",
      x"FFDD8E30",
      x"FFDD8627",
      x"FFD57D22",
      x"FFDA872C",
      x"FFDA8831",
      x"FFD88635",
      x"FFDD8C39",
      x"FFDF9138",
      x"FFDE9038",
      x"FFDF9335",
      x"FFDF9334",
      x"FFD88931",
      x"FFDC882D",
      x"FFE58625",
      x"FFE27B1B",
      x"FFE6801E",
      x"FFEE902D",
      x"FFEB8C29",
      x"FFEA8929",
      x"FFEF9330",
      x"FFE98D2B",
      x"FFE68427",
      x"FFE48222",
      x"FFE48324",
      x"FFE7872A",
      x"FFE88B2F",
      x"FFEA8E30",
      x"FFEB9035",
      x"FFED9841",
      x"FFED9A45",
      x"FFEA9542",
      x"FFE8913F",
      x"FFE68E3C",
      x"FFE9903D",
      x"FFE99241",
      x"FFE78C39",
      x"FFE48935",
      x"FFDC721C",
      x"FFE0751C",
      x"FFDC741E",
      x"FFE27F1D",
      x"FFEC9728",
      x"FFEC9225",
      x"FFF2A22F",
      x"FFEE9323",
      x"FFE57D16",
      x"FFE17510",
      x"FFE3831F",
      x"FFD87218",
      x"FFD47119",
      x"FFD16A19",
      x"FFD7771D",
      x"FFD36A12",
      x"FFD26F11",
      x"FFCF6D11",
      x"FFD06D11",
      x"FFE28921",
      x"FFE49833",
      x"FFD79236",
      x"FFD4872E",
      x"FFDB8A2B",
      x"FFDC8727",
      x"FFD77C23",
      x"FFD9862D",
      x"FFDA8A35",
      x"FFD88231",
      x"FFDC8A36",
      x"FFDF8E36",
      x"FFDD8F36",
      x"FFE09638",
      x"FFDE9034",
      x"FFD78229",
      x"FFDD8A2E",
      x"FFE98C2A",
      x"FFE27719",
      x"FFE88320",
      x"FFED902B",
      x"FFEB8C2A",
      x"FFE9892B",
      x"FFEF9432",
      x"FFEA8B29",
      x"FFE7882A",
      x"FFE68524",
      x"FFE07D20",
      x"FFE78729",
      x"FFEA8C2D",
      x"FFEA8C2C",
      x"FFE7903A",
      x"FFE78D35",
      x"FFEE9A44",
      x"FFEB943E",
      x"FFE78E3A",
      x"FFE38A3A",
      x"FFEA8E38",
      x"FFEA9546",
      x"FFEA8F3B",
      x"FFE48530",
      x"FFDC751F",
      x"FFE0761E",
      x"FFDC741F",
      x"FFDF771A",
      x"FFE89127",
      x"FFE8881E",
      x"FFF09C29",
      x"FFEF9426",
      x"FFE77E15",
      x"FFE47810",
      x"FFE5811A",
      x"FFDB771A",
      x"FFD06713",
      x"FFD36B19",
      x"FFD8771B",
      x"FFD67016",
      x"FFD37113",
      x"FFD16F13",
      x"FFD67211",
      x"FFE58D22",
      x"FFE59933",
      x"FFDA9439",
      x"FFD48832",
      x"FFDC8B2D",
      x"FFDF8827",
      x"FFD97D21",
      x"FFD68028",
      x"FFDA8932",
      x"FFDB8633",
      x"FFDC8834",
      x"FFDE8E37",
      x"FFDE9136",
      x"FFDD9033",
      x"FFDC8E33",
      x"FFD7842C",
      x"FFDD892D",
      x"FFEA8F2B",
      x"FFE58522",
      x"FFE7821C",
      x"FFEC8E2C",
      x"FFEB8D2A",
      x"FFEB8E2E",
      x"FFEC8E2C",
      x"FFEA8A27",
      x"FFE78729",
      x"FFE58424",
      x"FFE38020",
      x"FFE78728",
      x"FFE88C2D",
      x"FFEC902F",
      x"FFE48C38",
      x"FFE4882D",
      x"FFEE9C4A",
      x"FFED9945",
      x"FFE78D35",
      x"FFE58C3C",
      x"FFEB923C",
      x"FFEC9541",
      x"FFEA9242",
      x"FFE5842C",
      x"FFDE761F",
      x"FFE1761C",
      x"FFE07921",
      x"FFDD7419",
      x"FFE68B27",
      x"FFE47F18",
      x"FFEF9C2C",
      x"FFEF9A2A",
      x"FFE8841C",
      x"FFE47711",
      x"FFE27D17",
      x"FFDC781A",
      x"FFD36813",
      x"FFD36D1A",
      x"FFD9781C",
      x"FFD56F15",
      x"FFD67315",
      x"FFD16E12",
      x"FFD77513",
      x"FFE89225",
      x"FFE59A37",
      x"FFD99234",
      x"FFD3832C",
      x"FFDD8B2C",
      x"FFDE8726",
      x"FFD97E20",
      x"FFD9862D",
      x"FFDB8931",
      x"FFDB8735",
      x"FFDB8732",
      x"FFDF8E35",
      x"FFDD9137",
      x"FFDD8F33",
      x"FFD78B36",
      x"FFD98429",
      x"FFDD882C",
      x"FFEA922F",
      x"FFE68624",
      x"FFE9841E",
      x"FFEC912A",
      x"FFED9130",
      x"FFEA8B29",
      x"FFEC8D2B",
      x"FFEA8A28",
      x"FFEA8B2A",
      x"FFE98A2A",
      x"FFE27F20",
      x"FFE58222",
      x"FFE68425",
      x"FFEB8E2E",
      x"FFE68C38",
      x"FFE78C31",
      x"FFEE9944",
      x"FFEB9542",
      x"FFEA8E37",
      x"FFE58936",
      x"FFEA8F38",
      x"FFED9541",
      x"FFEB9542",
      x"FFE98B32",
      x"FFE17D25",
      x"FFE3791F",
      x"FFDF7B23",
      x"FFDD741A",
      x"FFE28623",
      x"FFE17515",
      x"FFEF9B2F",
      x"FFF2A338",
      x"FFE9851E",
      x"FFE37612",
      x"FFE17713",
      x"FFDD7618",
      x"FFD67017",
      x"FFD5701B",
      x"FFD9761B",
      x"FFD87518",
      x"FFD57113",
      x"FFD47415",
      x"FFDA7715",
      x"FFE99326",
      x"FFE79C35",
      x"FFD89034",
      x"FFD58730",
      x"FFDE8E30",
      x"FFDD8928",
      x"FFDA7E22",
      x"FFD98329",
      x"FFDB8833",
      x"FFD98531",
      x"FFDD8833",
      x"FFDE8C33",
      x"FFDE933B",
      x"FFDC903A",
      x"FFD78C37",
      x"FFDB872B",
      x"FFDE8D30",
      x"FFEB902B",
      x"FFE88927",
      x"FFEA8820",
      x"FFED9129",
      x"FFEC902F",
      x"FFEC8E2C",
      x"FFEC8B27",
      x"FFEB8A26",
      x"FFEA8C2A",
      x"FFEB8F2E",
      x"FFE48222",
      x"FFE78525",
      x"FFE88A2C",
      x"FFEB8D2D",
      x"FFE88C37",
      x"FFE98C31",
      x"FFED9844",
      x"FFED9644",
      x"FFE68D39",
      x"FFE68934",
      x"FFEA9038",
      x"FFEC9644",
      x"FFEC9340",
      x"FFEA9343",
      x"FFE2802C",
      x"FFE17820",
      x"FFDF7820",
      x"FFDC7016",
      x"FFDF7B1A",
      x"FFDE791A",
      x"FFED9A30",
      x"FFF0A339",
      x"FFEA8B22",
      x"FFE27610",
      x"FFE27710",
      x"FFDB7016",
      x"FFD6721A",
      x"FFD36B18",
      x"FFDA781D",
      x"FFD97518",
      x"FFD67515",
      x"FFD57315",
      x"FFDC7B14",
      x"FFE79224",
      x"FFE89C38",
      x"FFD78E30",
      x"FFD58833",
      x"FFDE8F30",
      x"FFDE8C2D",
      x"FFD87C21",
      x"FFD78227",
      x"FFDB842F",
      x"FFDA8332",
      x"FFDE8933",
      x"FFDD8A31",
      x"FFDC913B",
      x"FFD6862F",
      x"FFCF7F2B",
      x"FFDA8326",
      x"FFE28E2F",
      x"FFE68826",
      x"FFE88D2A",
      x"FFE88621",
      x"FFEA8924",
      x"FFE98C2A",
      x"FFEB8F2E",
      x"FFEC8D2C",
      x"FFEA8825",
      x"FFE98A28",
      x"FFE88929",
      x"FFE38421",
      x"FFE78926",
      x"FFE88B2C",
      x"FFEC912E",
      x"FFEA923A",
      x"FFE88B31",
      x"FFED9A46",
      x"FFEB9847",
      x"FFE58C3B",
      x"FFE48937",
      x"FFE88D38",
      x"FFED9643",
      x"FFEB9443",
      x"FFE89042",
      x"FFE1802C",
      x"FFDE731B",
      x"FFE27E25",
      x"FFDC7219",
      x"FFE2811E",
      x"FFDF781A",
      x"FFEA942D",
      x"FFF0A239",
      x"FFEC9127",
      x"FFE57C15",
      x"FFE37A13",
      x"FFDC7215",
      x"FFD7721B",
      x"FFD46C1A",
      x"FFDC7D21",
      x"FFD9771B",
      x"FFD57416",
      x"FFD57616",
      x"FFDD7B15",
      x"FFE89323",
      x"FFE69B37",
      x"FFD78D30",
      x"FFD6882F",
      x"FFE19134",
      x"FFDD8A2C",
      x"FFD77D22",
      x"FFD78127",
      x"FFDC8631",
      x"FFDB8633",
      x"FFDD8531",
      x"FFDE8C34",
      x"FFDD923B",
      x"FFD98C36",
      x"FFD27F2B",
      x"FFDA8226",
      x"FFE29134",
      x"FFE78926",
      x"FFE88D28",
      x"FFE47C1B",
      x"FFEA8B23",
      x"FFE98B28",
      x"FFEC8E2C",
      x"FFED8C2A",
      x"FFEB8B27",
      x"FFEB8D2B",
      x"FFE98928",
      x"FFE48322",
      x"FFE88726",
      x"FFE7892B",
      x"FFEC8E2B",
      x"FFEC953E",
      x"FFE68B32",
      x"FFEE9840",
      x"FFEB9746",
      x"FFE88E3B",
      x"FFE38838",
      x"FFE78A33",
      x"FFEB9445",
      x"FFEC9649",
      x"FFE99141",
      x"FFE38332",
      x"FFDE6E18",
      x"FFE27D23",
      x"FFDB7019",
      x"FFE1791A",
      x"FFDE791A",
      x"FFE98B25",
      x"FFF09D33",
      x"FFEC962E",
      x"FFE57C16",
      x"FFE07512",
      x"FFDA6D13",
      x"FFD56E19",
      x"FFD8721D",
      x"FFDA781C",
      x"FFD87419",
      x"FFD06F14",
      x"FFD47314",
      x"FFDB7713",
      x"FFE89324",
      x"FFE49A36",
      x"FFD89033",
      x"FFD78830",
      x"FFE19436",
      x"FFDD8C2D",
      x"FFD57C22",
      x"FFD37D26",
      x"FFDD8730",
      x"FFDC8533",
      x"FFDE8834",
      x"FFDF8D34",
      x"FFE0953F",
      x"FFDA9039",
      x"FFD47A26",
      x"FFDB8429",
      x"FFE28F33",
      x"FFE58725",
      x"FFE88B27",
      x"FFE68121",
      x"FFE6841F",
      x"FFEA8D2B",
      x"FFED9333",
      x"FFEE902D",
      x"FFE98828",
      x"FFEB8F2B",
      x"FFE88A2B",
      x"FFE38021",
      x"FFE98A29",
      x"FFE98A2C",
      x"FFEC912E",
      x"FFED9237",
      x"FFE88F36",
      x"FFEA923C",
      x"FFEB9747",
      x"FFE89140",
      x"FFE38A3D",
      x"FFE58734",
      x"FFEB9544",
      x"FFEC984A",
      x"FFE78D3C",
      x"FFE38738",
      x"FFDB6D18",
      x"FFE27C24",
      x"FFDA6D17",
      x"FFDD7419",
      x"FFDF791B",
      x"FFE68420",
      x"FFEF9B32",
      x"FFEE9930",
      x"FFE6821A",
      x"FFE17713",
      x"FFD86C14",
      x"FFD8751E",
      x"FFDA761D",
      x"FFDB791D",
      x"FFDA791A",
      x"FFD47317",
      x"FFD47515",
      x"FFD97714",
      x"FFE6962A",
      x"FFE09533",
      x"FFD89134",
      x"FFD8892F",
      x"FFE19535",
      x"FFDD8E2F",
      x"FFD17B22",
      x"FFD37E27",
      x"FFDA832D",
      x"FFDC8431",
      x"FFDB8330",
      x"FFDD8B31",
      x"FFDC8E35",
      x"FFDC913F",
      x"FFD77A21",
      x"FFDD872C",
      x"FFE39236",
      x"FFE28324",
      x"FFE88B26",
      x"FFE78622",
      x"FFE88720",
      x"FFEA8B27",
      x"FFE98D2B",
      x"FFEC8C2A",
      x"FFE98828",
      x"FFE88828",
      x"FFE78A2B",
      x"FFE07F23",
      x"FFE78A28",
      x"FFE88A2B",
      x"FFEB8E2F",
      x"FFEB9034",
      x"FFE98E35",
      x"FFEB933A",
      x"FFEB9B4A",
      x"FFE79242",
      x"FFE58E41",
      x"FFE48633",
      x"FFEA903B",
      x"FFED9849",
      x"FFEA9244",
      x"FFE48735",
      x"FFDA6B18",
      x"FFDD741D",
      x"FFD96E17",
      x"FFD97018",
      x"FFE07D1F",
      x"FFE4821E",
      x"FFEF9A33",
      x"FFEF9C34",
      x"FFE67B16",
      x"FFE17915",
      x"FFD96D13",
      x"FFD76F18",
      x"FFDB761C",
      x"FFDE7D20",
      x"FFDC7A1A",
      x"FFD57316",
      x"FFD37415",
      x"FFD97816",
      x"FFE49428",
      x"FFDB902F",
      x"FFD88E34",
      x"FFD88A30",
      x"FFE29738",
      x"FFDC8C2C",
      x"FFCA7820",
      x"FFD07D26",
      x"FFD7842E",
      x"FFDD8430",
      x"FFDC832F",
      x"FFDE8B33",
      x"FFDD9039",
      x"FFDB8E39",
      x"FFD77C22",
      x"FFDD892E",
      x"FFE29034",
      x"FFE08023",
      x"FFE58723",
      x"FFE6821E",
      x"FFE5821E",
      x"FFEB902C",
      x"FFE98927",
      x"FFE98C2B",
      x"FFEA8B28",
      x"FFE88B2A",
      x"FFE98B2C",
      x"FFE17E23",
      x"FFE68625",
      x"FFE88A2D",
      x"FFEB8E2F",
      x"FFEB9036",
      x"FFEC9238",
      x"FFEA923B",
      x"FFEF9D4B",
      x"FFE89140",
      x"FFE58D3E",
      x"FFE48634",
      x"FFEC9541",
      x"FFED9646",
      x"FFEB984D",
      x"FFE89241",
      x"FFDC6E1B",
      x"FFDD731C",
      x"FFDA721C",
      x"FFD86B13",
      x"FFDC781B",
      x"FFE3811D",
      x"FFEC9329",
      x"FFEF9E36",
      x"FFE98923",
      x"FFE27C17",
      x"FFDC7519",
      x"FFD8721A",
      x"FFDC791E",
      x"FFDE8023",
      x"FFDC7E1D",
      x"FFD67416",
      x"FFD27113",
      x"FFD77814",
      x"FFE49228",
      x"FFDC9131",
      x"FFD68B31",
      x"FFDD8D30",
      x"FFDC9135",
      x"FFD98A2D",
      x"FFCC7A21",
      x"FFCD7B25",
      x"FFD3802C",
      x"FFDD852F",
      x"FFDD8530",
      x"FFDD8A33",
      x"FFDC8F3A",
      x"FFDC8F3B",
      x"FFDC8429",
      x"FFE08B30",
      x"FFE29136",
      x"FFE38322",
      x"FFE58320",
      x"FFE47D1B",
      x"FFE4831F",
      x"FFE98F2A",
      x"FFE78728",
      x"FFEA8C2C",
      x"FFEB8F2D",
      x"FFEA8927",
      x"FFE8892A",
      x"FFE07D20",
      x"FFE58828",
      x"FFE88E30",
      x"FFEC9232",
      x"FFEB9033",
      x"FFEB9239",
      x"FFE88E37",
      x"FFED9A49",
      x"FFEA9544",
      x"FFE69044",
      x"FFE38534",
      x"FFEC9748",
      x"FFEF9D50",
      x"FFED994D",
      x"FFE58938",
      x"FFDD6F1D",
      x"FFDB6E1B",
      x"FFDA6F1B",
      x"FFD46613",
      x"FFD97218",
      x"FFE17D1D",
      x"FFE98D27",
      x"FFEF9D34",
      x"FFEB8D25",
      x"FFE27B18",
      x"FFDE781B",
      x"FFDA741E",
      x"FFDC781F",
      x"FFDC7D22",
      x"FFDE801E",
      x"FFD57415",
      x"FFD37416",
      x"FFDC7E18",
      x"FFE0902A",
      x"FFD98E33",
      x"FFD98C32",
      x"FFDE8E33",
      x"FFD78A30",
      x"FFD7892C",
      x"FFCC7C23",
      x"FFD08028",
      x"FFD07C29",
      x"FFD87F2C",
      x"FFDD8330",
      x"FFDE8B34",
      x"FFDA8C33",
      x"FFDB8D37",
      x"FFD98027",
      x"FFDF8A2F",
      x"FFE29338",
      x"FFE68724",
      x"FFE98A22",
      x"FFE37B1A",
      x"FFE47E1B",
      x"FFE78B27",
      x"FFE38524",
      x"FFE68829",
      x"FFEB8E2E",
      x"FFE98928",
      x"FFE98B2B",
      x"FFE17E22",
      x"FFE58627",
      x"FFE78A2C",
      x"FFEB8F2F",
      x"FFEB8C2D",
      x"FFEC933B",
      x"FFEA913B",
      x"FFEF9E4B",
      x"FFEA9340",
      x"FFE79042",
      x"FFE48A3D",
      x"FFED9543",
      x"FFEE9A4B",
      x"FFED9A50",
      x"FFE78E3E",
      x"FFDA6E1D",
      x"FFDA6E19",
      x"FFDB711C",
      x"FFD66412",
      x"FFDA7018",
      x"FFDF7818",
      x"FFE78A26",
      x"FFEE9A33",
      x"FFEB932A",
      x"FFE17B18",
      x"FFDC761A",
      x"FFDB7820",
      x"FFDD7B21",
      x"FFDD7F23",
      x"FFDC7C1B",
      x"FFD47315",
      x"FFD47416",
      x"FFD97A17",
      x"FFE08F28",
      x"FFDB9032",
      x"FFDC8F34",
      x"FFE29639",
      x"FFE39837",
      x"FFDA8C2E",
      x"FFD17D22",
      x"FFD18229",
      x"FFCE7B28",
      x"FFDA812E",
      x"FFDD822E",
      x"FFDD8931",
      x"FFDC8C33",
      x"FFD98934",
      x"FFD9822A",
      x"FFE08C32",
      x"FFE3963C",
      x"FFE38222",
      x"FFE27F1E",
      x"FFE57F1B",
      x"FFE17815",
      x"FFE78924",
      x"FFE68826",
      x"FFEA8B2A",
      x"FFEC8E2E",
      x"FFE88827",
      x"FFE98A2B",
      x"FFE17F24",
      x"FFE58527",
      x"FFE78B2D",
      x"FFE88B2E",
      x"FFEB8E30",
      x"FFEC9239",
      x"FFEA8F36",
      x"FFEF9D48",
      x"FFE9913D",
      x"FFE68D3F",
      x"FFE68E41",
      x"FFEA9441",
      x"FFEF9A4B",
      x"FFEE9D55",
      x"FFE78F40",
      x"FFD96B1C",
      x"FFDC6E1C",
      x"FFDB711B",
      x"FFD66814",
      x"FFD76B15",
      x"FFE07818",
      x"FFE37F1D",
      x"FFEB922C",
      x"FFEC942A",
      x"FFE17C18",
      x"FFDB7419",
      x"FFDB771F",
      x"FFDB761E",
      x"FFDF8224",
      x"FFDD7D1D",
      x"FFD37114",
      x"FFD47616",
      x"FFD97B18",
      x"FFE1912C",
      x"FFDD9237",
      x"FFDD9137",
      x"FFE49638",
      x"FFE49739",
      x"FFDA8E2F",
      x"FFD17D23",
      x"FFD2822A",
      x"FFCC7A28",
      x"FFD8802D",
      x"FFDE8430",
      x"FFDD872E",
      x"FFDC8B30",
      x"FFD88730",
      x"FFDE892E",
      x"FFE18E32",
      x"FFE4953A"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
