library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_white_queen_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_white_queen_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"40000000",
      x"82000000",
      x"82000000",
      x"40000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0D000000",
      x"45000000",
      x"5E000000",
      x"50000000",
      x"15000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"06000000",
      x"90000000",
      x"EE000000",
      x"FF000000",
      x"FF000000",
      x"EE000000",
      x"90000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0D000000",
      x"91000000",
      x"EA000000",
      x"F3000000",
      x"EE000000",
      x"D1000000",
      x"25000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"64000000",
      x"F9000000",
      x"FE262626",
      x"FFA8A8A8",
      x"FFA8A8A8",
      x"FE252525",
      x"F9000000",
      x"63000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"28000000",
      x"A6000000",
      x"C4000000",
      x"8E000000",
      x"19000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"60000000",
      x"FF000000",
      x"FE171717",
      x"FF363636",
      x"FF212121",
      x"FF030303",
      x"CF000000",
      x"15000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"BE000000",
      x"FF080808",
      x"FF888888",
      x"FFFAFAFA",
      x"FFFAFAFA",
      x"FF888888",
      x"FF080808",
      x"BC000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"51000000",
      x"FF000000",
      x"FF050505",
      x"FE0A0A0A",
      x"FF010101",
      x"C3000000",
      x"20000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"D9000000",
      x"FF141414",
      x"FFA9A9A9",
      x"FFF6F6F6",
      x"FFC7C7C7",
      x"FF212121",
      x"EE000000",
      x"50000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"B8000000",
      x"FF070707",
      x"FF828282",
      x"FFF9F9F9",
      x"FFF9F9F9",
      x"FF818181",
      x"FF070707",
      x"B7000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2E000000",
      x"DE000000",
      x"FF0C0C0C",
      x"FF646464",
      x"FF939393",
      x"FE4C4C4C",
      x"FF020202",
      x"8F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FD000000",
      x"FF2D2D2D",
      x"FFDEDEDE",
      x"FFFEFEFE",
      x"FFF7F7F7",
      x"FF363636",
      x"F3000000",
      x"5D000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"5F000000",
      x"FF000000",
      x"FF1A1A1A",
      x"FF757575",
      x"FF757575",
      x"FF1A1A1A",
      x"FF000000",
      x"5E000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"5A000000",
      x"F2000000",
      x"FF303030",
      x"FFE9E9E9",
      x"FFFCFCFC",
      x"FFCFCFCF",
      x"FF242424",
      x"F2000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0D000000",
      x"3D000000",
      x"7E000000",
      x"83000000",
      x"3C000000",
      x"0E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"BB000000",
      x"FF030303",
      x"FF929292",
      x"FFDBDBDB",
      x"FFA7A7A7",
      x"FE171717",
      x"E8000000",
      x"44000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"9E000000",
      x"F3000000",
      x"FE000000",
      x"FE000000",
      x"F3000000",
      x"9D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"59000000",
      x"F2000000",
      x"FF303030",
      x"FFE9E9E9",
      x"FFFBFBFB",
      x"FFCFCFCF",
      x"FF242424",
      x"F2000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"3C000000",
      x"83000000",
      x"7E000000",
      x"3D000000",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"16000000",
      x"95000000",
      x"F3000000",
      x"FE000000",
      x"FE000000",
      x"F5000000",
      x"88000000",
      x"0E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"41000000",
      x"E1000000",
      x"FF030303",
      x"FE292929",
      x"FE121212",
      x"FF000000",
      x"8F000000",
      x"0E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"89000000",
      x"F7000000",
      x"F7000000",
      x"89000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2E000000",
      x"DD000000",
      x"FE0B0B0B",
      x"FF626262",
      x"FF8F8F8F",
      x"FF4C4C4C",
      x"FF010101",
      x"8E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"89000000",
      x"F5000000",
      x"FE000000",
      x"FE000000",
      x"F3000000",
      x"95000000",
      x"16000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"61000000",
      x"F1000000",
      x"FE161616",
      x"FF9C9C9C",
      x"FFAEAEAE",
      x"FE0E0E0E",
      x"F5000000",
      x"3B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"04000000",
      x"3F000000",
      x"C9000000",
      x"FF000000",
      x"ED000000",
      x"66000000",
      x"0E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"6C000000",
      x"F5000000",
      x"F5000000",
      x"6C000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"50000000",
      x"FF000000",
      x"FE040404",
      x"FE090909",
      x"FF010101",
      x"C2000000",
      x"20000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3C000000",
      x"F5000000",
      x"FE0F0F0F",
      x"FFAEAEAE",
      x"FF9C9C9C",
      x"FE161616",
      x"F1000000",
      x"60000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"8F000000",
      x"FB000000",
      x"FF6D6D6D",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFACACAC",
      x"FF000000",
      x"7F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"65000000",
      x"FF000000",
      x"F5000000",
      x"41000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"8D000000",
      x"FB000000",
      x"FB000000",
      x"8D000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3B000000",
      x"EE000000",
      x"FF000000",
      x"AB000000",
      x"18000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"80000000",
      x"FF000000",
      x"FFADADAD",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FF6C6C6C",
      x"FB000000",
      x"8F000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"8E000000",
      x"FB000000",
      x"FF6F6F6F",
      x"FFFDFDFD",
      x"FFFEFEFE",
      x"FF9B9B9B",
      x"FF000000",
      x"7B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF000000",
      x"FE000000",
      x"AA000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"AB000000",
      x"FF000000",
      x"FF000000",
      x"AB000000",
      x"0F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"66000000",
      x"FC000000",
      x"FF000000",
      x"65000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"7C000000",
      x"FF000000",
      x"FF9B9B9B",
      x"FFFEFEFE",
      x"FFFDFDFD",
      x"FF6E6E6E",
      x"FB000000",
      x"8E000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"60000000",
      x"F3000000",
      x"FE131313",
      x"FF6E6E6E",
      x"FF6D6D6D",
      x"FE151515",
      x"F5000000",
      x"3E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF000000",
      x"FF000000",
      x"F9000000",
      x"27000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1D000000",
      x"C8000000",
      x"FE010101",
      x"FE010101",
      x"C8000000",
      x"1D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"E3000000",
      x"FF000000",
      x"FF000000",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3E000000",
      x"F5000000",
      x"FE161616",
      x"FF6D6D6D",
      x"FF6E6E6E",
      x"FE131313",
      x"F3000000",
      x"60000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"A8000000",
      x"F3000000",
      x"FB000000",
      x"FE000000",
      x"FF000000",
      x"AC000000",
      x"0F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF000000",
      x"FF010101",
      x"FF000000",
      x"9B000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2D000000",
      x"E7000000",
      x"FF2F2F2F",
      x"FF2F2F2F",
      x"E7000000",
      x"2D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"5D000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"AB000000",
      x"FF000000",
      x"FE000000",
      x"FB000000",
      x"F3000000",
      x"A8000000",
      x"0F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"12000000",
      x"5E000000",
      x"8B000000",
      x"D3000000",
      x"FF000000",
      x"CF000000",
      x"24000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF141414",
      x"FE060606",
      x"DA000000",
      x"25000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"45000000",
      x"FD000000",
      x"FF707070",
      x"FF707070",
      x"FD000000",
      x"45000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"10000000",
      x"C2000000",
      x"FF010101",
      x"FF060606",
      x"FF010101",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"25000000",
      x"CF000000",
      x"FE000000",
      x"D2000000",
      x"8B000000",
      x"5E000000",
      x"12000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"08000000",
      x"79000000",
      x"FF000000",
      x"FD000000",
      x"A6000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF030303",
      x"FF494949",
      x"FF1F1F1F",
      x"F1000000",
      x"5E000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"7B000000",
      x"FF000000",
      x"FFB0B0B0",
      x"FFB0B0B0",
      x"FF000000",
      x"7B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"46000000",
      x"EA000000",
      x"FF121212",
      x"FF2F2F2F",
      x"FF030303",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"A6000000",
      x"FD000000",
      x"FF000000",
      x"79000000",
      x"08000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"3C000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"5B000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF6C6C6C",
      x"FF656565",
      x"FC000000",
      x"9D000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"C0000000",
      x"FF0D0D0D",
      x"FFCBCBCB",
      x"FFCBCBCB",
      x"FF0D0D0D",
      x"C0000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"07000000",
      x"84000000",
      x"F9000000",
      x"FF3F3F3F",
      x"FF626262",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"5B000000",
      x"FF000000",
      x"FE000000",
      x"FF000000",
      x"3C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"DA000000",
      x"2C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF666666",
      x"FFD6D6D6",
      x"FE0B0B0B",
      x"D7000000",
      x"23000000",
      x"00000000",
      x"00000000",
      x"06000000",
      x"F5000000",
      x"FF2C2C2C",
      x"FFDCDCDC",
      x"FFDCDCDC",
      x"FF2C2C2C",
      x"F5000000",
      x"06000000",
      x"00000000",
      x"00000000",
      x"1A000000",
      x"C2000000",
      x"FF000000",
      x"FFB2B2B2",
      x"FF696969",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2C000000",
      x"D9000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"DE000000",
      x"FF101010",
      x"FF0B0B0B",
      x"FB000000",
      x"8F000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FF666666",
      x"FC000000",
      x"5E000000",
      x"00000000",
      x"00000000",
      x"35000000",
      x"FF000000",
      x"FF4B4B4B",
      x"FFECECEC",
      x"FFECECEC",
      x"FF4B4B4B",
      x"FF000000",
      x"35000000",
      x"00000000",
      x"00000000",
      x"40000000",
      x"F8000000",
      x"FF3B3B3B",
      x"FFF1F1F1",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"8F000000",
      x"FB000000",
      x"FF0B0B0B",
      x"FF101010",
      x"DE000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"A5000000",
      x"FF090909",
      x"FF8E8E8E",
      x"FE0D0D0D",
      x"E6000000",
      x"3B000000",
      x"00000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFC8C8C8",
      x"FF090909",
      x"D3000000",
      x"04000000",
      x"00000000",
      x"79000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"79000000",
      x"00000000",
      x"01000000",
      x"B2000000",
      x"FF050505",
      x"FFB2B2B2",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"00000000",
      x"3B000000",
      x"E5000000",
      x"FE0D0D0D",
      x"FF8E8E8E",
      x"FF090909",
      x"A5000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"6C000000",
      x"FF000000",
      x"FFA9A9A9",
      x"FF898989",
      x"FE080808",
      x"C3000000",
      x"13000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFE8E8E8",
      x"FE434343",
      x"FF000000",
      x"4E000000",
      x"00000000",
      x"B4000000",
      x"FF080808",
      x"FF868686",
      x"FFFAFAFA",
      x"FFFAFAFA",
      x"FF868686",
      x"FF080808",
      x"B4000000",
      x"00000000",
      x"33000000",
      x"FD000000",
      x"FF333333",
      x"FFE1E1E1",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"13000000",
      x"C3000000",
      x"FE080808",
      x"FF8A8A8A",
      x"FFA9A9A9",
      x"FF000000",
      x"6C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"40000000",
      x"FF000000",
      x"FF6D6D6D",
      x"FFE9E9E9",
      x"FE464646",
      x"FE000000",
      x"98000000",
      x"00000000",
      x"68000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFF9F9F9",
      x"FF808080",
      x"FF070707",
      x"B9000000",
      x"17000000",
      x"CE000000",
      x"FE0D0D0D",
      x"FFA6A6A6",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFA6A6A6",
      x"FE0D0D0D",
      x"CE000000",
      x"13000000",
      x"AB000000",
      x"FF040404",
      x"FF707070",
      x"FFF5F5F5",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"68000000",
      x"00000000",
      x"98000000",
      x"FE000000",
      x"FF464646",
      x"FFE9E9E9",
      x"FF6D6D6D",
      x"FF000000",
      x"40000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2F000000",
      x"EB000000",
      x"FF333333",
      x"FFFDFDFD",
      x"FFAAAAAA",
      x"FE111111",
      x"E9000000",
      x"48000000",
      x"69000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFBBBBBB",
      x"FF151515",
      x"E2000000",
      x"66000000",
      x"DE000000",
      x"FF191919",
      x"FFC2C2C2",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFC2C2C2",
      x"FF191919",
      x"DE000000",
      x"5B000000",
      x"DD000000",
      x"FE121212",
      x"FFB1B1B1",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"69000000",
      x"48000000",
      x"E9000000",
      x"FE111111",
      x"FFA9A9A9",
      x"FFFDFDFD",
      x"FF333333",
      x"EB000000",
      x"2F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"21000000",
      x"D1000000",
      x"FF070707",
      x"FFFBFBFB",
      x"FFF1F1F1",
      x"FF606060",
      x"FD000000",
      x"A5000000",
      x"78000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFF0F0F0",
      x"FF3D3D3D",
      x"F6000000",
      x"C1000000",
      x"F2000000",
      x"FF2A2A2A",
      x"FFE1E1E1",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE1E1E1",
      x"FF2A2A2A",
      x"F2000000",
      x"B9000000",
      x"F4000000",
      x"FF343434",
      x"FFEAEAEA",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"78000000",
      x"A5000000",
      x"FC000000",
      x"FF606060",
      x"FFF1F1F1",
      x"FFFBFBFB",
      x"FF070707",
      x"D1000000",
      x"22000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"B7000000",
      x"FE000000",
      x"FFD5D5D5",
      x"FFFFFFFF",
      x"FFEDEDED",
      x"FE1E1E1E",
      x"F5000000",
      x"C1000000",
      x"FF020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF9E9E9E",
      x"FE000000",
      x"FA000000",
      x"FE000000",
      x"FF3A3A3A",
      x"FFFCFCFC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFCFCFC",
      x"FF3A3A3A",
      x"FE000000",
      x"F9000000",
      x"FE000000",
      x"FF8E8E8E",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FF020202",
      x"C1000000",
      x"F5000000",
      x"FE1E1E1E",
      x"FFEDEDED",
      x"FFFFFFFF",
      x"FFD5D5D5",
      x"FE000000",
      x"B7000000",
      x"13000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"A1000000",
      x"FE000000",
      x"FF9B9B9B",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFBBBBBB",
      x"FE0A0A0A",
      x"FF000000",
      x"FE020202",
      x"FF656565",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF151515",
      x"FF000000",
      x"FF000000",
      x"FF6E6E6E",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF6E6E6E",
      x"FF000000",
      x"FF000000",
      x"FF0F0F0F",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF4F4F4",
      x"FF656565",
      x"FE020202",
      x"FF000000",
      x"FE0B0B0B",
      x"FFBBBBBB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF9B9B9B",
      x"FE000000",
      x"A1000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"07000000",
      x"86000000",
      x"FA000000",
      x"FF636363",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFF1F1F1",
      x"FF636363",
      x"FF040404",
      x"FF020202",
      x"FF676767",
      x"FFF5F5F5",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF888888",
      x"FF000000",
      x"FF000000",
      x"FF999999",
      x"FFE0E0E0",
      x"FFDEDEDE",
      x"FFDDDDDD",
      x"FFDFDFDF",
      x"FF979797",
      x"FF000000",
      x"FF000000",
      x"FF7A7A7A",
      x"FFF4F4F4",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFF5F5F5",
      x"FF686868",
      x"FF020202",
      x"FF040404",
      x"FF656565",
      x"FFF0F0F0",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FF626262",
      x"FA000000",
      x"86000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"6B000000",
      x"F5000000",
      x"FF3E3E3E",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFBDBDBD",
      x"FF191919",
      x"FF010101",
      x"FF313131",
      x"FF606060",
      x"FF4A4A4A",
      x"FF3F3F3F",
      x"FF3B3B3B",
      x"FF282828",
      x"FF000000",
      x"FF000000",
      x"FF212121",
      x"FF2A2A2A",
      x"FF282828",
      x"FF282828",
      x"FF292929",
      x"FF202020",
      x"FF000000",
      x"FF000000",
      x"FF232323",
      x"FF353535",
      x"FF3A3A3A",
      x"FF3D3D3D",
      x"FF464646",
      x"FF212121",
      x"FF000000",
      x"FF121212",
      x"FFA4A4A4",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF3E3E3E",
      x"F5000000",
      x"6B000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"53000000",
      x"F0000000",
      x"FF171717",
      x"FF646464",
      x"FF3F3F3F",
      x"FF0A0A0A",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF020202",
      x"FF040404",
      x"FF070707",
      x"FF090909",
      x"FF0B0B0B",
      x"FF0C0C0C",
      x"FF0D0D0D",
      x"FF0E0E0E",
      x"FF0F0F0F",
      x"FF101010",
      x"FF111111",
      x"FF111111",
      x"FF101010",
      x"FF0F0F0F",
      x"FF0E0E0E",
      x"FF0D0D0D",
      x"FF0C0C0C",
      x"FF0B0B0B",
      x"FF090909",
      x"FF070707",
      x"FF040404",
      x"FF020202",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF202020",
      x"FF535353",
      x"FF141414",
      x"F0000000",
      x"53000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"41000000",
      x"E8000000",
      x"FF000000",
      x"FF000000",
      x"FF0A0A0A",
      x"FF202020",
      x"FF343434",
      x"FF474747",
      x"FF575757",
      x"FF646464",
      x"FF747474",
      x"FF818181",
      x"FF8D8D8D",
      x"FF989898",
      x"FFA0A0A0",
      x"FFA7A7A7",
      x"FFAAAAAA",
      x"FFADADAD",
      x"FFB0B0B0",
      x"FFB1B1B1",
      x"FFB1B1B1",
      x"FFB0B0B0",
      x"FFADADAD",
      x"FFAAAAAA",
      x"FFA7A7A7",
      x"FFA0A0A0",
      x"FF989898",
      x"FF8D8D8D",
      x"FF818181",
      x"FF747474",
      x"FF646464",
      x"FF575757",
      x"FF474747",
      x"FF343434",
      x"FF202020",
      x"FF0A0A0A",
      x"FF000000",
      x"FF000000",
      x"E6000000",
      x"3F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"28000000",
      x"D9000000",
      x"FF0A0A0A",
      x"FF828282",
      x"FFCACACA",
      x"FFD5D5D5",
      x"FFE0E0E0",
      x"FFEBEBEB",
      x"FFF1F1F1",
      x"FFF4F4F4",
      x"FFF7F7F7",
      x"FFF9F9F9",
      x"FFFBFBFB",
      x"FFFDFDFD",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFDFDFD",
      x"FFFBFBFB",
      x"FFF9F9F9",
      x"FFF7F7F7",
      x"FFF4F4F4",
      x"FFF1F1F1",
      x"FFEBEBEB",
      x"FFE0E0E0",
      x"FFD5D5D5",
      x"FFCACACA",
      x"FF818181",
      x"FF0A0A0A",
      x"D9000000",
      x"27000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"B1000000",
      x"FF030303",
      x"FE5A5A5A",
      x"FFE7E7E7",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFE7E7E7",
      x"FF5A5A5A",
      x"FF030303",
      x"B1000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2C000000",
      x"CA000000",
      x"FF070707",
      x"FE5C5C5C",
      x"FFECECEC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFECECEC",
      x"FF5B5B5B",
      x"FF060606",
      x"CA000000",
      x"2C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"30000000",
      x"CC000000",
      x"FF030303",
      x"FF5F5F5F",
      x"FFFCFCFC",
      x"FFEEEEEE",
      x"FFC9C9C9",
      x"FFA8A8A8",
      x"FF8D8D8D",
      x"FF767676",
      x"FF686868",
      x"FF575757",
      x"FF494949",
      x"FF3D3D3D",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3B3B3B",
      x"FF3D3D3D",
      x"FF494949",
      x"FF585858",
      x"FF686868",
      x"FF767676",
      x"FF8E8E8E",
      x"FFA8A8A8",
      x"FFC9C9C9",
      x"FFEEEEEE",
      x"FFFCFCFC",
      x"FF5E5E5E",
      x"FF030303",
      x"CB000000",
      x"2F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"4A000000",
      x"EA000000",
      x"FE020202",
      x"FF0A0A0A",
      x"FF0C0C0C",
      x"FF111111",
      x"FF171717",
      x"FF1C1C1C",
      x"FF232323",
      x"FF272727",
      x"FF2C2C2C",
      x"FF303030",
      x"FF343434",
      x"FF363636",
      x"FF373737",
      x"FF383838",
      x"FF393939",
      x"FF393939",
      x"FF383838",
      x"FF373737",
      x"FF363636",
      x"FF343434",
      x"FF303030",
      x"FF2C2C2C",
      x"FF272727",
      x"FF232323",
      x"FF1C1C1C",
      x"FF161616",
      x"FF111111",
      x"FF0C0C0C",
      x"FF0A0A0A",
      x"FE020202",
      x"E9000000",
      x"49000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"8B000000",
      x"FF000000",
      x"FE1A1A1A",
      x"FF929292",
      x"FFB3B3B3",
      x"FFC2C2C2",
      x"FFCFCFCF",
      x"FFD9D9D9",
      x"FFE0E0E0",
      x"FFE7E7E7",
      x"FFEEEEEE",
      x"FFF4F4F4",
      x"FFF7F7F7",
      x"FFF9F9F9",
      x"FFFAFAFA",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFAFAFA",
      x"FFF9F9F9",
      x"FFF6F6F6",
      x"FFF4F4F4",
      x"FFEEEEEE",
      x"FFE7E7E7",
      x"FFE0E0E0",
      x"FFD9D9D9",
      x"FFCFCFCF",
      x"FFC2C2C2",
      x"FFB4B4B4",
      x"FF909090",
      x"FE1A1A1A",
      x"FF000000",
      x"8C000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0D000000",
      x"C1000000",
      x"FF060606",
      x"FFC6C6C6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFC6C6C6",
      x"FF060606",
      x"C1000000",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"84000000",
      x"FF010101",
      x"FFBFBFBF",
      x"FFFDFDFD",
      x"FFF9F9F9",
      x"FFF7F7F7",
      x"FFF4F4F4",
      x"FFF2F2F2",
      x"FFF0F0F0",
      x"FFEDEDED",
      x"FFE9E9E9",
      x"FFE6E6E6",
      x"FFE3E3E3",
      x"FFE2E2E2",
      x"FFE1E1E1",
      x"FFE1E1E1",
      x"FFE2E2E2",
      x"FFE3E3E3",
      x"FFE6E6E6",
      x"FFE9E9E9",
      x"FFEDEDED",
      x"FFF0F0F0",
      x"FFF2F2F2",
      x"FFF4F4F4",
      x"FFF7F7F7",
      x"FFF9F9F9",
      x"FFFDFDFD",
      x"FFBEBEBE",
      x"FF010101",
      x"83000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"C8000000",
      x"FF050505",
      x"FF868686",
      x"FF979797",
      x"FF828282",
      x"FF727272",
      x"FF626262",
      x"FF595959",
      x"FF535353",
      x"FF4C4C4C",
      x"FF444444",
      x"FF3E3E3E",
      x"FF3A3A3A",
      x"FF383838",
      x"FF343434",
      x"FF343434",
      x"FF383838",
      x"FF3A3A3A",
      x"FF3E3E3E",
      x"FF444444",
      x"FF4C4C4C",
      x"FF535353",
      x"FF595959",
      x"FF626262",
      x"FF727272",
      x"FF828282",
      x"FF979797",
      x"FF878787",
      x"FF050505",
      x"C8000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"79000000",
      x"FB000000",
      x"FF010101",
      x"FF0B0B0B",
      x"FF0E0E0E",
      x"FF272727",
      x"FF454545",
      x"FF626262",
      x"FF7E7E7E",
      x"FF939393",
      x"FFA5A5A5",
      x"FFB7B7B7",
      x"FFC2C2C2",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC2C2C2",
      x"FFB7B7B7",
      x"FFA5A5A5",
      x"FF939393",
      x"FF7E7E7E",
      x"FF626262",
      x"FF454545",
      x"FF272727",
      x"FF0E0E0E",
      x"FF0B0B0B",
      x"FF010101",
      x"FB000000",
      x"70000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"4B000000",
      x"EB000000",
      x"FE0B0B0B",
      x"FF6A6A6A",
      x"FFD7D7D7",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFBFBFB",
      x"FFFAFAFA",
      x"FFF9F9F9",
      x"FFF7F7F7",
      x"FFF6F6F6",
      x"FFF5F5F5",
      x"FFF5F5F5",
      x"FFF5F5F5",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF4F4F4",
      x"FFF5F5F5",
      x"FFF5F5F5",
      x"FFF6F6F6",
      x"FFF7F7F7",
      x"FFF8F8F8",
      x"FFF9F9F9",
      x"FFFBFBFB",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD7D7D7",
      x"FF676767",
      x"FE080808",
      x"E2000000",
      x"34000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0B000000",
      x"97000000",
      x"FC000000",
      x"FF444444",
      x"FFB7B7B7",
      x"FFB3B3B3",
      x"FFA8A8A8",
      x"FF9E9E9E",
      x"FF909090",
      x"FF858585",
      x"FF7D7D7D",
      x"FF757575",
      x"FF6E6E6E",
      x"FF686868",
      x"FF666666",
      x"FF636363",
      x"FF616161",
      x"FF606060",
      x"FF606060",
      x"FF626262",
      x"FF656565",
      x"FF676767",
      x"FF6C6C6C",
      x"FF737373",
      x"FF7B7B7B",
      x"FF838383",
      x"FF8C8C8C",
      x"FF999999",
      x"FFA5A5A5",
      x"FFAFAFAF",
      x"FFBDBDBD",
      x"FFBFBFBF",
      x"FF2A2A2A",
      x"F4000000",
      x"63000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"21000000",
      x"D1000000",
      x"FE000000",
      x"FF101010",
      x"FF181818",
      x"FF111111",
      x"FF0E0E0E",
      x"FF0C0C0C",
      x"FF141414",
      x"FF232323",
      x"FF313131",
      x"FF3E3E3E",
      x"FF4B4B4B",
      x"FF555555",
      x"FF5C5C5C",
      x"FF5E5E5E",
      x"FF626262",
      x"FF676767",
      x"FF626262",
      x"FF5F5F5F",
      x"FF5D5D5D",
      x"FF565656",
      x"FF515151",
      x"FF434343",
      x"FF363636",
      x"FF282828",
      x"FF1A1A1A",
      x"FF0B0B0B",
      x"FF0D0D0D",
      x"FF101010",
      x"FF151515",
      x"FF1E1E1E",
      x"FF090909",
      x"F8000000",
      x"7B000000",
      x"06000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"64000000",
      x"FF000000",
      x"FF292929",
      x"FF787878",
      x"FFA5A5A5",
      x"FFCACACA",
      x"FFE5E5E5",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF0F0F0",
      x"FFD3D3D3",
      x"FFB3B3B3",
      x"FF888888",
      x"FF414141",
      x"FF020202",
      x"BB000000",
      x"15000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"9E000000",
      x"FE000000",
      x"FFA0A0A0",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF0F0F0",
      x"FF161616",
      x"E3000000",
      x"2B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"5C000000",
      x"FF000000",
      x"FE1E1E1E",
      x"FF474747",
      x"FF727272",
      x"FF9D9D9D",
      x"FFC4C4C4",
      x"FFE1E1E1",
      x"FFFCFCFC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFCFCFC",
      x"FFE1E1E1",
      x"FFC4C4C4",
      x"FF9C9C9C",
      x"FF727272",
      x"FF474747",
      x"FE060606",
      x"D4000000",
      x"23000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"12000000",
      x"A4000000",
      x"F1000000",
      x"F7000000",
      x"FA000000",
      x"FE000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF060606",
      x"FF1C1C1C",
      x"FF2D2D2D",
      x"FF3D3D3D",
      x"FF4C4C4C",
      x"FF585858",
      x"FF5D5D5D",
      x"FF626262",
      x"FF696969",
      x"FF696969",
      x"FF626262",
      x"FF5D5D5D",
      x"FF585858",
      x"FF4C4C4C",
      x"FF3D3D3D",
      x"FF2D2D2D",
      x"FF1C1C1C",
      x"FF060606",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FE000000",
      x"FA000000",
      x"F7000000",
      x"EF000000",
      x"85000000",
      x"09000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1B000000",
      x"5A000000",
      x"76000000",
      x"8B000000",
      x"A0000000",
      x"AC000000",
      x"B8000000",
      x"C5000000",
      x"D1000000",
      x"DA000000",
      x"E2000000",
      x"E9000000",
      x"F0000000",
      x"F4000000",
      x"F6000000",
      x"F9000000",
      x"FB000000",
      x"FB000000",
      x"F9000000",
      x"F6000000",
      x"F4000000",
      x"F0000000",
      x"E9000000",
      x"E2000000",
      x"DA000000",
      x"D1000000",
      x"C5000000",
      x"B8000000",
      x"AC000000",
      x"A0000000",
      x"8B000000",
      x"76000000",
      x"59000000",
      x"17000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"05000000",
      x"08000000",
      x"0C000000",
      x"0F000000",
      x"14000000",
      x"1B000000",
      x"22000000",
      x"26000000",
      x"2B000000",
      x"2E000000",
      x"32000000",
      x"34000000",
      x"35000000",
      x"37000000",
      x"38000000",
      x"38000000",
      x"37000000",
      x"35000000",
      x"34000000",
      x"32000000",
      x"2E000000",
      x"2B000000",
      x"26000000",
      x"22000000",
      x"1B000000",
      x"14000000",
      x"0F000000",
      x"0C000000",
      x"08000000",
      x"05000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
