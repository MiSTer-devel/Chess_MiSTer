library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_black_mister_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_black_mister_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF282827",
      x"FFA7A6A6",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB7B7B6",
      x"FF3E3E3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF6A6A6A",
      x"FF0F0E0E",
      x"FF272727",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF302F2F",
      x"FF080807",
      x"FF8B8A8A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA8A7A7",
      x"FF292828",
      x"FFEBEBEB",
      x"FF9B9B9B",
      x"FF373737",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF50504F",
      x"FF8F8F8F",
      x"FFECECEC",
      x"FF383737",
      x"FFC7C6C6",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF373636",
      x"FF8F8E8E",
      x"FFFFFFFF",
      x"FFFBFBFB",
      x"FF515150",
      x"FF6D6D6D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF939392",
      x"FF50504F",
      x"FFF9F8F8",
      x"FFFFFFFF",
      x"FF8B8B8B",
      x"FF676666",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA3A2A2",
      x"FF3D3D3D",
      x"FFE6E6E5",
      x"00000000",
      x"FF98CAAD",
      x"FFD8D8D7",
      x"FF2F2F2E",
      x"FFABABAA",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF292929",
      x"FFD2D2D2",
      x"FF9BCCB0",
      x"00000000",
      x"FFE3E4E4",
      x"FF3B3B3B",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464545",
      x"FF8B8A89",
      x"FFF6FBF8",
      x"00000000",
      x"00000000",
      x"FFF8FCFA",
      x"FF9E9E9D",
      x"FF313131",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF4F4F4E",
      x"FF959595",
      x"FFF9FCFA",
      x"00000000",
      x"00000000",
      x"FFF4FAF8",
      x"FF848483",
      x"FF6B6B6A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF9D9D9D",
      x"FF0A0A09",
      x"FFE7E7E7",
      x"FFF4F4F4",
      x"FFE8E8E8",
      x"FFE7E6E7",
      x"FFEFEFEF",
      x"FFF3F3F3",
      x"FF2C2B2A",
      x"FF535252",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF7B7C7B",
      x"FF232222",
      x"FFF2F2F2",
      x"FFEFEFEF",
      x"FFE7E7E7",
      x"FFE8E8E8",
      x"FFF4F4F4",
      x"FFECECEC",
      x"FF212121",
      x"FFC9C9C9",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF373635",
      x"FF0E0D0C",
      x"FF504F4E",
      x"FF555454",
      x"FF3E3E3E",
      x"FF3D3C3D",
      x"FF4C4B4A",
      x"FF545352",
      x"FF181716",
      x"FF0B0A09",
      x"FF797877",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF8C8B8A",
      x"FF878686",
      x"FF181716",
      x"FF161514",
      x"FF535252",
      x"FF4C4B4A",
      x"FF3D3D3D",
      x"FF3E3E3E",
      x"FF545353",
      x"FF515050",
      x"FF0D0C0C",
      x"FF7C7C7C",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF505050",
      x"FF0C0C0C",
      x"FF11100F",
      x"FF1A1918",
      x"FF121110",
      x"FF121110",
      x"FF161514",
      x"FF171615",
      x"FF131211",
      x"FF121110",
      x"FF191817",
      x"FF1A1918",
      x"FF090907",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF181716",
      x"FF191817",
      x"FF121110",
      x"FF131211",
      x"FF171514",
      x"FF161514",
      x"FF121110",
      x"FF121110",
      x"FF181716",
      x"FF121111",
      x"FF474646",
      x"FFA1A1A1",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF595858",
      x"FF0D0C0B",
      x"FF161514",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF161514",
      x"FF11100F",
      x"FF121211",
      x"FF8B8A8A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF8C8C8B",
      x"FF0A0909",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF141413",
      x"FFADADAC",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF4E4E4D",
      x"FF11100F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF0F0F0E",
      x"FF626262",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF424241",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF3D3C3C",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF454444",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF3D3D3C",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464645",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF3D3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464645",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF3D3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464645",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF141312",
      x"FF171616",
      x"FF171616",
      x"FF141312",
      x"FF181716",
      x"FF181716",
      x"FF141312",
      x"FF181717",
      x"FF161615",
      x"FF151313",
      x"FF191716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF3D3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464645",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF141312",
      x"FF1E1E1D",
      x"FFBBBABA",
      x"FFBDBCBC",
      x"FF201F1E",
      x"FF141312",
      x"FF141312",
      x"FF242423",
      x"FFC1C0C0",
      x"FFB6B6B6",
      x"FF1A1A19",
      x"FF151413",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF3D3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464645",
      x"FF0B0B0A",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF100F0D",
      x"FF0B0A09",
      x"FF6A6A69",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF7B7A7A",
      x"FF0D0C0B",
      x"FF0A0A09",
      x"FF7C7C7C",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF616060",
      x"FF0A0909",
      x"FF0F0E0D",
      x"FF0F0E0D",
      x"FF0F0E0D",
      x"FF0F0E0D",
      x"FF0F0E0E",
      x"FF100F0E",
      x"FF0F0E0D",
      x"FF0F0E0D",
      x"FF100F0E",
      x"FF100F0D",
      x"FF0F0E0D",
      x"FF100F0E",
      x"FF100F0E",
      x"FF100F0D",
      x"FF0B0B0A",
      x"FF3D3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF464645",
      x"FF494948",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA5A5A5",
      x"FFA2A2A1",
      x"FFC1C0C0",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFDEDEDE",
      x"FF979797",
      x"FF8E8E8E",
      x"FFD7D6D6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFB8B7B7",
      x"FF979797",
      x"FF9C9C9B",
      x"FF9C9C9B",
      x"FF9E9D9C",
      x"FF9E9D9C",
      x"FF9F9E9E",
      x"FF9F9F9E",
      x"FFA1A09F",
      x"FFA1A0A0",
      x"FFA2A1A1",
      x"FFA2A2A2",
      x"FFA3A3A3",
      x"FFA4A3A3",
      x"FFA5A4A4",
      x"FFA5A5A5",
      x"FF444443",
      x"FF3E3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF3C3B3B",
      x"FFA4A4A4",
      x"FFFEFEFE",
      x"FFFAFAFA",
      x"FFF9F9F9",
      x"FFF9F9F9",
      x"FFF9F9F9",
      x"FFF9F9F9",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFBFBFB",
      x"FFF9F9F9",
      x"FFF9F9F9",
      x"FFF9F9F9",
      x"FFFAFAFA",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFDFDFD",
      x"FFFDFDFD",
      x"FFFCFCFC",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFCFCFC",
      x"FFFAFAFA",
      x"FFFAFAFA",
      x"FFFAFAFA",
      x"FFFAFAFA",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FF9F9F9E",
      x"FF363635",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF3A3939",
      x"FFB2B1B1",
      x"FFF0F0F0",
      x"FF7F7F7F",
      x"FF555555",
      x"FF555555",
      x"FF555555",
      x"FF555555",
      x"FF878787",
      x"FFF9F9F9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF818181",
      x"FF555555",
      x"FF555555",
      x"FF555555",
      x"FF656565",
      x"FFD6D6D6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD9D9D9",
      x"FF717171",
      x"FF616161",
      x"FF616161",
      x"FF606060",
      x"FF8E8E8E",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF6F6F6",
      x"FF898989",
      x"FF595959",
      x"FF585858",
      x"FF575757",
      x"FF565656",
      x"FF808080",
      x"FFF3F3F3",
      x"FFAFAFAF",
      x"FF333332",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF383737",
      x"FFACABAB",
      x"FFEFEFEF",
      x"FF464646",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF323232",
      x"FFDCDCDC",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFEEEEEE",
      x"FF141414",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF181818",
      x"FFC2C2C2",
      x"FFF0F0F0",
      x"FF9F9F9C",
      x"FFA4A4A1",
      x"FFF3F3F2",
      x"FFBCBCBC",
      x"FF121212",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF181818",
      x"FFF1F1F1",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD8D8D8",
      x"FF2E2E2E",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF4B4B4B",
      x"FFF4F4F4",
      x"FFA9A9A9",
      x"FF333333",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF434342",
      x"FF949394",
      x"FFFDFDFD",
      x"FF6C6C6C",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF070707",
      x"FF676767",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFEBEBEB",
      x"FF696969",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF333333",
      x"FFDDDDDD",
      x"FFE0E0DF",
      x"FF6B6A66",
      x"FF6C6B68",
      x"FFE2E2E1",
      x"FFD8D8D8",
      x"FF2E2E2E",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF707070",
      x"FFEDEDED",
      x"FFFFFFFF",
      x"FFF2F2F2",
      x"FF616161",
      x"FF060606",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF777777",
      x"FFFEFEFE",
      x"FF8E8D8D",
      x"FF3C3C3B",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA6A5A5",
      x"FF201F1F",
      x"FF50504F",
      x"FFFFFFFF",
      x"FFD4D4D4",
      x"FF040404",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF131313",
      x"FF343434",
      x"FF111111",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF787878",
      x"FFFEFEFE",
      x"FFEDEDEC",
      x"FFCECECD",
      x"FFD0D0CF",
      x"FFF0F0F0",
      x"FFFCFCFC",
      x"FF717171",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF131313",
      x"FF333333",
      x"FF111111",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF070707",
      x"FFDADADA",
      x"FFFFFFFF",
      x"FF494847",
      x"FF100F0F",
      x"FF757575",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF383838",
      x"FF111010",
      x"FF121110",
      x"FF121211",
      x"FFE2E2E2",
      x"FFFFFFFF",
      x"FF565656",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF323232",
      x"FFE6E6E6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE4E4E4",
      x"FF656565",
      x"FF0D0D0D",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF5F5F5F",
      x"FFFEFEFE",
      x"FFDCDCDB",
      x"FF11100F",
      x"FF141312",
      x"FF10100F",
      x"FF2F2F2F",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC6C6C6",
      x"FF252525",
      x"FF11100F",
      x"FF191817",
      x"FF181716",
      x"FF0E0D0C",
      x"FF5D5D5C",
      x"FFF1F1F1",
      x"FFE3E3E3",
      x"FF555555",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF0A0A0A",
      x"FF8A8A8A",
      x"FFF0F0F0",
      x"FFE9E9E9",
      x"FFFDFEFD",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFF4FBF7",
      x"FFE4E4E3",
      x"FFE9E9E9",
      x"FFCBCBCB",
      x"FF272727",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF5A5A5A",
      x"FFE6E6E6",
      x"FFF0F0F0",
      x"FF575757",
      x"FF100F0E",
      x"FF181716",
      x"FF191817",
      x"FF11100F",
      x"FF282727",
      x"FFCBCACA",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF545353",
      x"FF0D0D0C",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF161615",
      x"FF929291",
      x"FFFFFFFF",
      x"FFE2E2E2",
      x"FF555555",
      x"FF070707",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF070707",
      x"FF7E7E7E",
      x"FFF5F5F5",
      x"FFA2A1A1",
      x"FF6E6D6C",
      x"FFF4F4F4",
      x"FFDEF1E8",
      x"00000000",
      x"00000000",
      x"FFDCF0E6",
      x"FFFAFBFB",
      x"FF81817F",
      x"FF5F5F5D",
      x"FFE2E2E1",
      x"FFBDBDBD",
      x"FF262626",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF090909",
      x"FF5A5A5A",
      x"FFE4E4E4",
      x"FFFFFFFF",
      x"FF8B8B8B",
      x"FF151514",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF0D0C0C",
      x"FF565555",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF060606",
      x"FF161514",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF161514",
      x"FF070706",
      x"FF909090",
      x"FFF0F0F0",
      x"FFFEFEFE",
      x"FFC9C9C9",
      x"FF646464",
      x"FF3A3A3A",
      x"FF282828",
      x"FF262626",
      x"FF333333",
      x"FF4C4C4C",
      x"FFACACAC",
      x"FFF8F8F8",
      x"FF999998",
      x"FF363633",
      x"FF3E3D3B",
      x"FF403F3E",
      x"FFB4B4B4",
      x"FFF7F6F6",
      x"FFF8F7F8",
      x"FFBABAB9",
      x"FF464543",
      x"FF3F3E3C",
      x"FF393836",
      x"FF5E5D5B",
      x"FFEEEEEE",
      x"FFC1C1C1",
      x"FF4A4A4A",
      x"FF323232",
      x"FF262626",
      x"FF282828",
      x"FF3B3B3B",
      x"FF666666",
      x"FFCDCDCD",
      x"FFFFFFFF",
      x"FFEFEFEF",
      x"FF8B8A8A",
      x"FF090908",
      x"FF171615",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF171615",
      x"FF070606",
      x"FFC9C9C9",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF9F9F9E",
      x"FF080808",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF161514",
      x"FF141313",
      x"FF5F5F5F",
      x"FFDFDFDF",
      x"FFFFFFFF",
      x"FFFAFAFA",
      x"FFE4E4E4",
      x"FFD2D2D2",
      x"FFD0D0D0",
      x"FFDDDDDD",
      x"FFF2F2F2",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFD0D0D0",
      x"FF5B5A58",
      x"FF3F3E3C",
      x"FF373634",
      x"FF4A4947",
      x"FF6D6B6A",
      x"FF6F6E6C",
      x"FF4E4D4B",
      x"FF363533",
      x"FF42413F",
      x"FF3F3E3C",
      x"FFB1B0AF",
      x"FFF7F7F7",
      x"FFFFFFFF",
      x"FFF1F1F1",
      x"FFDCDCDC",
      x"FFD0D0D0",
      x"FFD2D2D2",
      x"FFE5E5E5",
      x"FFFAFAFA",
      x"FFFFFFFF",
      x"FFDCDCDC",
      x"FF5C5C5C",
      x"FF141413",
      x"FF171514",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF090808",
      x"FF8B8B8A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF868685",
      x"FF080807",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF0E0D0D",
      x"FF131312",
      x"FF545454",
      x"FFA8A9A9",
      x"FFC8C8C8",
      x"FFD6D6D6",
      x"FFD8D8D8",
      x"FFCFCFCF",
      x"FFF5F5F5",
      x"FFFFFFFF",
      x"FF9E9E9D",
      x"FF3A3939",
      x"FF7D7C7B",
      x"FF383735",
      x"FF3A3937",
      x"FF343331",
      x"FF81807F",
      x"FF848483",
      x"FF31302E",
      x"FF3E3D3B",
      x"FF3A3937",
      x"FF696867",
      x"FF585755",
      x"FF6C6C6A",
      x"FFF4F4F4",
      x"FFFDFCFC",
      x"FFDADADA",
      x"FFD6D6D6",
      x"FFD6D6D6",
      x"FFC8C7C7",
      x"FFA7A7A7",
      x"FF525150",
      x"FF131212",
      x"FF0E0D0D",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF0A0908",
      x"FF6E6E6D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF888888",
      x"FF080807",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF151413",
      x"FF100F0F",
      x"FF111110",
      x"FF1E1E1E",
      x"FF2C2C2C",
      x"FF2E2E2E",
      x"FF5D5D5D",
      x"FFB6B6B6",
      x"FFC8C7C7",
      x"FFD4D4D3",
      x"FFC5C4C4",
      x"FF797876",
      x"FF272624",
      x"FF484746",
      x"FFA8A8A7",
      x"FFF1F1F1",
      x"FFEFEFEF",
      x"FF91908F",
      x"FF3C3B39",
      x"FF2A2926",
      x"FF545351",
      x"FFCCCCCC",
      x"FFD4D4D4",
      x"FFD7D7D7",
      x"FF9E9E9D",
      x"FF9F9F9F",
      x"FF2C2C2C",
      x"FF2C2C2C",
      x"FF1E1D1D",
      x"FF111010",
      x"FF100F0F",
      x"FF151413",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF090808",
      x"FF717170",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB3B3B2",
      x"FF080807",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF141312",
      x"FF141312",
      x"FFDADADA",
      x"FF3E3E3E",
      x"FF595959",
      x"FFEEEEEE",
      x"FFF0F0F0",
      x"FFCBCACA",
      x"FFE0DFDF",
      x"FFF6F6F6",
      x"FFE0E0DF",
      x"FFE1E1E0",
      x"FFE2E2E1",
      x"FFE8E8E7",
      x"FFF5F5F4",
      x"FFD8D8D7",
      x"FFD3D3D2",
      x"FFF0F0F0",
      x"FFE8E8E8",
      x"FF8B8B8B",
      x"FF1A1A1A",
      x"FFC2C2C1",
      x"FF474646",
      x"FF111010",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF090808",
      x"FF999999",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF1C1B1B",
      x"FF141312",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF5F5E5E",
      x"FFB1B0B0",
      x"FF090909",
      x"FFBEBEBE",
      x"FF7D7D7D",
      x"FF7E7D7D",
      x"FFBBBBBA",
      x"FFFFFFFF",
      x"FFF1F1F1",
      x"FF9C9B98",
      x"FF888885",
      x"FF888783",
      x"FFA2A29F",
      x"FFF5F5F5",
      x"FFFFFFFF",
      x"FFC7C7C7",
      x"FF797878",
      x"FF545353",
      x"FFC6C6C6",
      x"FF181717",
      x"FF717171",
      x"FFA5A4A4",
      x"FF0F0E0E",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF141312",
      x"FF0C0C0C",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA5A5A5",
      x"FF161514",
      x"FF161514",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF0D0D0C",
      x"FFA4A4A3",
      x"FF757575",
      x"FF383837",
      x"FFBFBFBE",
      x"FF181716",
      x"FF090807",
      x"FF060605",
      x"FF727171",
      x"FFC4C4C4",
      x"FFEBEBEB",
      x"FFFBFBFB",
      x"FFFCFCFC",
      x"FFEEEEEE",
      x"FFCCCCCC",
      x"FF828282",
      x"FF0B0A0A",
      x"FF0A0908",
      x"FF0B0B0A",
      x"FF929292",
      x"FF8D8D8D",
      x"FF1E1D1C",
      x"FFC9C9C9",
      x"FF20201F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF171615",
      x"FF141413",
      x"FF8D8D8C",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF8E8E8E",
      x"FF040404",
      x"FF121110",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF0F0E0E",
      x"FF7E7D7D",
      x"FF50504F",
      x"FF818080",
      x"FF9A9999",
      x"FF0E0D0D",
      x"FF181716",
      x"FF161514",
      x"FF10100E",
      x"FF1E1E1E",
      x"FF454545",
      x"FF656564",
      x"FF686767",
      x"FF494949",
      x"FF222222",
      x"FF100F0F",
      x"FF151413",
      x"FF181716",
      x"FF11100F",
      x"FF4B4A4A",
      x"FFB4B3B3",
      x"FF131312",
      x"FF9B9A99",
      x"FF21201F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF141312",
      x"FF070606",
      x"FF747474",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBFBEBE",
      x"FF535353",
      x"FF161514",
      x"FF171615",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF0E0D0C",
      x"FF040404",
      x"FFA3A3A3",
      x"FF7A7A7A",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF151412",
      x"FF0E0D0C",
      x"FF0D0C0B",
      x"FF131211",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF282726",
      x"FFC7C7C6",
      x"FF1D1D1D",
      x"FF0B0A09",
      x"FF171615",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF151414",
      x"FF444444",
      x"FFA5A5A4",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF41413F",
      x"FF111010",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF121110",
      x"FF5C5B5A",
      x"FF4B4A4A",
      x"FF141312",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF141413",
      x"FF20201F",
      x"FF6F6E6D",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF111110",
      x"FF3E3D3D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF444342",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF0E0E0D",
      x"FF0F0E0D",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF171615",
      x"FF0C0C0B",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF454444",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF444342",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF444343",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF444342",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF444343",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF444342",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF444343",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF444342",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF454444",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF4A4948",
      x"FF100F0F",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF100F0F",
      x"FF474646",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBEBEBD",
      x"FF858585",
      x"FF252524",
      x"FF151413",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF121110",
      x"FF0E0E0D",
      x"FF0E0D0C",
      x"FF0E0D0C",
      x"FF0E0E0D",
      x"FF111010",
      x"FF171615",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF171615",
      x"FF191817",
      x"FF5A5A5A",
      x"FFB5B5B5",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB8B8B7",
      x"FF1C1C1B",
      x"FF0D0C0B",
      x"FF161514",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191716",
      x"FF171514",
      x"FF0A0909",
      x"FF2B2B2B",
      x"FF6D6D6C",
      x"FF888888",
      x"FF888888",
      x"FF6E6E6E",
      x"FF2E2D2C",
      x"FF0B0A09",
      x"FF161514",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF161514",
      x"FF0F0E0E",
      x"FF1B1B1B",
      x"FFB3B2B2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF3D3D3D",
      x"FF151413",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF100E0E",
      x"FF262626",
      x"FFAFAFAF",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB3B3B2",
      x"FF292928",
      x"FF0F0E0D",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181615",
      x"FF2E2D2D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF2F2E2E",
      x"FF191817",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF151413",
      x"FF292929",
      x"FFBEBEBE",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC2C2C2",
      x"FF2B2B2B",
      x"FF141312",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF191817",
      x"FF171616",
      x"FFC0BFBF",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF454544",
      x"FF131212",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF161514",
      x"FF100F0F",
      x"FFCACACA",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF111111",
      x"FF151413",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF181716",
      x"FF242424",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA9A7A8",
      x"FF030303",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF060606",
      x"FF535353",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF5A5A5A",
      x"FF050505",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF080807",
      x"FF070707",
      x"FF747473",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB4B4B4",
      x"FF7B7B7B",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7B7A79",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF7B7A7A",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7F7E7E",
      x"FF7D7C7B",
      x"FFA5A4A4",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
