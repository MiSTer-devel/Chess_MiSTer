library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_white_knight_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_white_knight_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"38000000",
      x"11000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"A1000000",
      x"98000000",
      x"13000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"14000000",
      x"C9000000",
      x"FF000000",
      x"DA000000",
      x"44000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"1F000000",
      x"C7000000",
      x"FF000000",
      x"FE000000",
      x"87000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"37000000",
      x"E2000000",
      x"FF020202",
      x"FF030303",
      x"E3000000",
      x"51000000",
      x"00000000",
      x"00000000",
      x"12000000",
      x"A5000000",
      x"FB000000",
      x"FE262626",
      x"FF191919",
      x"F0000000",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"39000000",
      x"E3000000",
      x"FF181818",
      x"FE505050",
      x"FE080808",
      x"DA000000",
      x"35000000",
      x"00000000",
      x"69000000",
      x"F8000000",
      x"FE272727",
      x"FFD2D2D2",
      x"FF4D4D4D",
      x"FF000000",
      x"2F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"2E000000",
      x"DD000000",
      x"FF1A1A1A",
      x"FFAFAFAF",
      x"FF424242",
      x"FC000000",
      x"CB000000",
      x"99000000",
      x"F7000000",
      x"FF111111",
      x"FFC9C9C9",
      x"FFF2F2F2",
      x"FF5B5B5B",
      x"FF000000",
      x"94000000",
      x"41000000",
      x"30000000",
      x"1E000000",
      x"0E000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0C000000",
      x"BF000000",
      x"FF080808",
      x"FF888888",
      x"FFCACACA",
      x"FF242424",
      x"FF000000",
      x"FF000000",
      x"FF050505",
      x"FF6A6A6A",
      x"FFF2F2F2",
      x"FFF7F7F7",
      x"FF7A7A7A",
      x"FF060606",
      x"FF000000",
      x"FE000000",
      x"EC000000",
      x"CB000000",
      x"A4000000",
      x"75000000",
      x"40000000",
      x"0C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"A5000000",
      x"FF040404",
      x"FF737373",
      x"FFF6F6F6",
      x"FFD8D8D8",
      x"FFC3C3C3",
      x"FFC3C3C3",
      x"FFC7C7C7",
      x"FFE7E7E7",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFE8E8E8",
      x"FCC6C6C6",
      x"FFA8A8A8",
      x"FF727272",
      x"FF313131",
      x"FE000000",
      x"FE000000",
      x"F7000000",
      x"E7000000",
      x"B7000000",
      x"33000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"22000000",
      x"D7000000",
      x"FE0D0D0D",
      x"FF9F9F9F",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FEFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF2F2F2",
      x"FF959595",
      x"FF414141",
      x"FE1B1B1B",
      x"FE060606",
      x"FF000000",
      x"99000000",
      x"23000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"83000000",
      x"F7000000",
      x"FF323232",
      x"FFE0E0E0",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF8F8F8",
      x"FFC4C4C4",
      x"FF7D7D7D",
      x"FE292929",
      x"FD000000",
      x"D0000000",
      x"62000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"48000000",
      x"EF000000",
      x"FE000000",
      x"FFC2C2C2",
      x"FFFBFBFB",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF8F8F8",
      x"FFDCDCDC",
      x"FF686868",
      x"FE000000",
      x"F2000000",
      x"93000000",
      x"07000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1A000000",
      x"FF000000",
      x"FF090909",
      x"FF959595",
      x"FFD8D8D8",
      x"FF3A3A3A",
      x"FF000000",
      x"FFC6C6C6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF6F6F6",
      x"FF818181",
      x"FE0D0D0D",
      x"F7000000",
      x"81000000",
      x"0A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"10000000",
      x"AE000000",
      x"FF030303",
      x"FF5F5F5F",
      x"FFDDDDDD",
      x"FF3C3C3C",
      x"FF000000",
      x"FF000000",
      x"FF787878",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF1F1F1",
      x"FF8A8A8A",
      x"FF050505",
      x"EB000000",
      x"6B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"56000000",
      x"EE000000",
      x"FE191919",
      x"FFBEBEBE",
      x"FF787878",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FFC3C3C3",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF8F8F8",
      x"FF868686",
      x"FF000000",
      x"F2000000",
      x"52000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"B1000000",
      x"FE000000",
      x"FF666666",
      x"FFF6F6F6",
      x"FF333333",
      x"FF000000",
      x"FF020202",
      x"FF444444",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFE8E8E8",
      x"FF464646",
      x"FE010101",
      x"DB000000",
      x"25000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"57000000",
      x"F2000000",
      x"FF2E2E2E",
      x"FFE9E9E9",
      x"FFF5F5F5",
      x"FF4D4D4D",
      x"FF030303",
      x"FF3D3D3D",
      x"FFD6D6D6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FFE6E6E6",
      x"FFEDEDED",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FFA7A7A7",
      x"FF111111",
      x"F9000000",
      x"87000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"06000000",
      x"E6000000",
      x"FF0A0A0A",
      x"FFB4B4B4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE0E0E0",
      x"FFC3C3C3",
      x"FFDFDFDF",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFECECEC",
      x"FF5C5C5C",
      x"FF3C3C3C",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF6F6F6",
      x"FF414141",
      x"FE000000",
      x"DD000000",
      x"26000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"04000000",
      x"92000000",
      x"FF010101",
      x"FF535353",
      x"FFEDEDED",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE0E0E0",
      x"FF333333",
      x"FF030303",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFC4C4C4",
      x"FF050505",
      x"FE000000",
      x"82000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"38000000",
      x"E3000000",
      x"FE111111",
      x"FFA8A8A8",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFC5C5C5",
      x"FF121212",
      x"FF313131",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FF575757",
      x"FE000000",
      x"F0000000",
      x"1F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"8C000000",
      x"FB000000",
      x"FF3E3E3E",
      x"FFF5F5F5",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FF474747",
      x"FF000000",
      x"FF9D9D9D",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFC0C0C0",
      x"FE0C0C0C",
      x"FF000000",
      x"94000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"29000000",
      x"D8000000",
      x"FE080808",
      x"FFC6C6C6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF9F9F9",
      x"FF8C8C8C",
      x"FF000000",
      x"FF272727",
      x"FFDADADA",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE6E6E6",
      x"FF3F3F3F",
      x"FE000000",
      x"D3000000",
      x"1A000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"8D000000",
      x"FF000000",
      x"FF6F6F6F",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFAFAFA",
      x"FFA6A6A6",
      x"FF141414",
      x"FF000000",
      x"FF343434",
      x"FFE0E0E0",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF6F6F6",
      x"FF717171",
      x"FF040404",
      x"EB000000",
      x"4B000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"29000000",
      x"F6000000",
      x"FF242424",
      x"FFD4D4D4",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFC5C5C5",
      x"FF1C1C1C",
      x"FF010101",
      x"FE000000",
      x"FF353535",
      x"FFE1E1E1",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFA3A3A3",
      x"FF0D0D0D",
      x"F7000000",
      x"79000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"06000000",
      x"B0000000",
      x"FF030303",
      x"FF6A6A6A",
      x"FFF5F5F5",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFF8F8F8",
      x"FFB9B9B9",
      x"FE050505",
      x"F7000000",
      x"9E000000",
      x"FF000000",
      x"FF3C3C3C",
      x"FFE5E5E5",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFCBCBCB",
      x"FF1E1E1E",
      x"FE000000",
      x"A5000000",
      x"0E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"39000000",
      x"E4000000",
      x"FF161616",
      x"FFB5B5B5",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF5F5F5",
      x"FF8F8F8F",
      x"FE131313",
      x"F6000000",
      x"8C000000",
      x"37000000",
      x"FF000000",
      x"FF4B4B4B",
      x"FFEDEDED",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF1F1F1",
      x"FF333333",
      x"FE000000",
      x"C7000000",
      x"1C000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"05000000",
      x"77000000",
      x"F7000000",
      x"FF3A3A3A",
      x"FFD4D4D4",
      x"FF585858",
      x"FF585858",
      x"FFDCDCDC",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF616161",
      x"FE0C0C0C",
      x"FF000000",
      x"7D000000",
      x"0D000000",
      x"5A000000",
      x"FF010101",
      x"FF5E5E5E",
      x"FFF3F3F3",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF585858",
      x"FF000000",
      x"EB000000",
      x"30000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"AA000000",
      x"FF000000",
      x"FF9B9B9B",
      x"FF7E7E7E",
      x"FF050505",
      x"FF050505",
      x"FF7A7A7A",
      x"FFF8F8F8",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFCFCFC",
      x"FFD5D5D5",
      x"FF3B3B3B",
      x"FE000000",
      x"E9000000",
      x"64000000",
      x"00000000",
      x"01000000",
      x"A0000000",
      x"FF060606",
      x"FF808080",
      x"FFF9F9F9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF9B9B9B",
      x"FF000000",
      x"FF000000",
      x"47000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1A000000",
      x"C3000000",
      x"FF000000",
      x"FFEDEDED",
      x"FF808080",
      x"FF060606",
      x"FF070707",
      x"FF808080",
      x"FFF8F8F8",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFFEFEFE",
      x"FFF4F4F4",
      x"FF9A9A9A",
      x"FE2E2E2E",
      x"FE020202",
      x"C6000000",
      x"4E000000",
      x"05000000",
      x"00000000",
      x"19000000",
      x"D2000000",
      x"FE0E0E0E",
      x"FFA6A6A6",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD8D8D8",
      x"FF000000",
      x"FF000000",
      x"82000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1B000000",
      x"C5000000",
      x"FF000000",
      x"FFFDFDFD",
      x"FFE7E7E7",
      x"FF8B8B8B",
      x"FF8B8B8B",
      x"FFE6E6E6",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE0E0E0",
      x"FF515151",
      x"FE0C0C0C",
      x"FF000000",
      x"96000000",
      x"1C000000",
      x"03000000",
      x"00000000",
      x"00000000",
      x"51000000",
      x"EE000000",
      x"FF232323",
      x"FFD4D4D4",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFCFCFC",
      x"FF030303",
      x"FF000000",
      x"BB000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"B6000000",
      x"FF000000",
      x"FFD8D8D8",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFDFDFD",
      x"FFC8C8C8",
      x"FF737373",
      x"FFA1A1A1",
      x"FFF3F3F3",
      x"FFFFFFFF",
      x"FFDEDEDE",
      x"FF484848",
      x"FF010101",
      x"E5000000",
      x"73000000",
      x"08000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0D000000",
      x"9D000000",
      x"FC000000",
      x"FF5B5B5B",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF2E2E2E",
      x"FF000000",
      x"EE000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0B000000",
      x"99000000",
      x"FD000000",
      x"FF818181",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFEEEEEE",
      x"FF4F4F4F",
      x"FF000000",
      x"FF121212",
      x"FFB4B4B4",
      x"FFE4E4E4",
      x"FF4B4B4B",
      x"FE000000",
      x"BE000000",
      x"44000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"4A000000",
      x"E8000000",
      x"FE1B1B1B",
      x"FFDBDBDB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF585858",
      x"FF000000",
      x"FF000000",
      x"0D000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"02000000",
      x"66000000",
      x"F4000000",
      x"FF202020",
      x"FFC3C3C3",
      x"FFFFFFFF",
      x"FFEAEAEA",
      x"FF434343",
      x"FF000000",
      x"FF191919",
      x"FFB9B9B9",
      x"FF545454",
      x"FF010101",
      x"BD000000",
      x"24000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1C000000",
      x"E5000000",
      x"FF030303",
      x"FFA3A3A3",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF7F7F7F",
      x"FF000000",
      x"FF000000",
      x"32000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1B000000",
      x"BC000000",
      x"FA000000",
      x"FF000000",
      x"FF111111",
      x"FF0B0B0B",
      x"FF000000",
      x"FF000000",
      x"FF3A3A3A",
      x"FF888888",
      x"FE0B0B0B",
      x"E1000000",
      x"3F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"21000000",
      x"D0000000",
      x"FF030303",
      x"FF5E5E5E",
      x"FFF0F0F0",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF9E9E9E",
      x"FF000000",
      x"FF000000",
      x"55000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"28000000",
      x"8C000000",
      x"C3000000",
      x"D7000000",
      x"D6000000",
      x"EB000000",
      x"FE000000",
      x"FE252525",
      x"FE1C1C1C",
      x"F2000000",
      x"60000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"20000000",
      x"AF000000",
      x"FB000000",
      x"FF3D3D3D",
      x"FFD4D4D4",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFB8B8B8",
      x"FF000000",
      x"FF000000",
      x"75000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"09000000",
      x"1A000000",
      x"25000000",
      x"25000000",
      x"7C000000",
      x"F6000000",
      x"FF010101",
      x"EE000000",
      x"5C000000",
      x"04000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0F000000",
      x"CC000000",
      x"FB000000",
      x"FE2C2C2C",
      x"FFE2E2E2",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFEFEFE",
      x"FFC3C3C3",
      x"FF000000",
      x"FF000000",
      x"8F000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"07000000",
      x"54000000",
      x"66000000",
      x"22000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"20000000",
      x"CC000000",
      x"FF020202",
      x"FF363636",
      x"FFE0E0E0",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFC7C7C7",
      x"FF060606",
      x"FF000000",
      x"A7000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"13000000",
      x"A7000000",
      x"FB000000",
      x"FF383838",
      x"FFC8C8C8",
      x"FFFDFDFD",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCACACA",
      x"FF0C0C0C",
      x"FF000000",
      x"B8000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"8D000000",
      x"F9000000",
      x"FE2B2B2B",
      x"FFE1E1E1",
      x"FFFDFDFD",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCDCDCD",
      x"FF111111",
      x"FF000000",
      x"C2000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"51000000",
      x"FF000000",
      x"FE202020",
      x"FFD5D5D5",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCFCFCF",
      x"FF141414",
      x"FF000000",
      x"C4000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1D000000",
      x"CF000000",
      x"FF090909",
      x"FF898989",
      x"FFF9F9F9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCFCFCF",
      x"FF141414",
      x"FF000000",
      x"C5000000",
      x"02000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"01000000",
      x"57000000",
      x"F0000000",
      x"FF262626",
      x"FFDADADA",
      x"FFFEFEFE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCFCFCF",
      x"FF141414",
      x"FF000000",
      x"C6000000",
      x"04000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"08000000",
      x"88000000",
      x"FA000000",
      x"FF5E5E5E",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCECECE",
      x"FF121212",
      x"FF000000",
      x"C7000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"0E000000",
      x"A9000000",
      x"FE000000",
      x"FFB7B7B7",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCCCCCC",
      x"FF0F0F0F",
      x"FF000000",
      x"C7000000",
      x"06000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"17000000",
      x"BD000000",
      x"FE000000",
      x"FFF4F4F4",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFD1D1D1",
      x"FF0A0A0A",
      x"FF000000",
      x"C7000000",
      x"05000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"1D000000",
      x"C8000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"C6000000",
      x"01000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"18000000",
      x"A2000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"CA000000",
      x"9E000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"03000000",
      x"18000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"1D000000",
      x"17000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
