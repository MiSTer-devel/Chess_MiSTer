library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_tile_0 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_tile_0 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"FF853301",
      x"FF833101",
      x"FF843203",
      x"FF863402",
      x"FF863402",
      x"FF863402",
      x"FF853301",
      x"FF8C3A02",
      x"FF8C3A02",
      x"FF8A3A02",
      x"FF8B3B01",
      x"FF8B3B02",
      x"FF883701",
      x"FF903E01",
      x"FF974402",
      x"FF924100",
      x"FF934202",
      x"FF8E3E02",
      x"FF8A3902",
      x"FF873702",
      x"FF8B3C02",
      x"FF934303",
      x"FF954501",
      x"FF974402",
      x"FF974402",
      x"FF944000",
      x"FF954101",
      x"FF954102",
      x"FF964302",
      x"FF944001",
      x"FF954201",
      x"FF9B4802",
      x"FF994601",
      x"FF9C4902",
      x"FF9D4B02",
      x"FF9B4901",
      x"FF9C4A01",
      x"FF9F4D03",
      x"FF9F4D03",
      x"FF9A4801",
      x"FF8A3902",
      x"FF8C3D03",
      x"FF8C3D02",
      x"FF8F4002",
      x"FF8C3D04",
      x"FF8D3E03",
      x"FF853702",
      x"FF8B3C04",
      x"FF873802",
      x"FF883902",
      x"FF893A02",
      x"FF873A01",
      x"FF883D02",
      x"FF863A01",
      x"FF8B3C02",
      x"FF8B3C01",
      x"FF8A3B02",
      x"FF883900",
      x"FF873800",
      x"FF863A01",
      x"FF863402",
      x"FF823000",
      x"FF812F01",
      x"FF853302",
      x"FF843201",
      x"FF853301",
      x"FF853302",
      x"FF893702",
      x"FF8D3B01",
      x"FF893801",
      x"FF8D3D01",
      x"FF883701",
      x"FF883603",
      x"FF8E3B00",
      x"FF964301",
      x"FF914001",
      x"FF924102",
      x"FF8C3C02",
      x"FF8A3902",
      x"FF853501",
      x"FF8A3A02",
      x"FF904002",
      x"FF954402",
      x"FF964301",
      x"FF964301",
      x"FF944001",
      x"FF933F00",
      x"FF933F02",
      x"FF954101",
      x"FF923E00",
      x"FF954201",
      x"FF994601",
      x"FF994601",
      x"FF9A4700",
      x"FF9D4B01",
      x"FF9B4802",
      x"FF9B4800",
      x"FF9D4B02",
      x"FF9D4B02",
      x"FF984601",
      x"FF873400",
      x"FF883901",
      x"FF8C3D03",
      x"FF8C3E01",
      x"FF893C02",
      x"FF893D02",
      x"FF823601",
      x"FF893C03",
      x"FF843702",
      x"FF823500",
      x"FF853800",
      x"FF8A3C03",
      x"FF873B00",
      x"FF853901",
      x"FF8B3E03",
      x"FF8D3E03",
      x"FF8A3B02",
      x"FF8A3B02",
      x"FF873800",
      x"FF893D02",
      x"FF863403",
      x"FF843201",
      x"FF823000",
      x"FF833102",
      x"FF853304",
      x"FF823001",
      x"FF833102",
      x"FF853301",
      x"FF8D3C05",
      x"FF883600",
      x"FF8C3A02",
      x"FF873501",
      x"FF863402",
      x"FF893601",
      x"FF934203",
      x"FF923E01",
      x"FF933F01",
      x"FF8E3A02",
      x"FF883602",
      x"FF843401",
      x"FF883701",
      x"FF8F3E02",
      x"FF923F01",
      x"FF934201",
      x"FF934201",
      x"FF914001",
      x"FF8F3E01",
      x"FF933F01",
      x"FF943E02",
      x"FF923C00",
      x"FF933F01",
      x"FF994403",
      x"FF994401",
      x"FF9B4701",
      x"FF9E4A02",
      x"FF9D4B03",
      x"FF994700",
      x"FF9C4A01",
      x"FF9C4A01",
      x"FF994502",
      x"FF893802",
      x"FF863A01",
      x"FF8A3C00",
      x"FF8D3E03",
      x"FF893902",
      x"FF883901",
      x"FF833601",
      x"FF893A05",
      x"FF863601",
      x"FF853502",
      x"FF853502",
      x"FF893A03",
      x"FF883803",
      x"FF863600",
      x"FF8A3B03",
      x"FF883901",
      x"FF8A3B02",
      x"FF863702",
      x"FF833701",
      x"FF833602",
      x"FF843202",
      x"FF843201",
      x"FF823001",
      x"FF812F01",
      x"FF823001",
      x"FF823001",
      x"FF833102",
      x"FF833101",
      x"FF8A3902",
      x"FF883501",
      x"FF8A3801",
      x"FF873600",
      x"FF863403",
      x"FF863301",
      x"FF913F04",
      x"FF903C01",
      x"FF923E01",
      x"FF8E3A01",
      x"FF883602",
      x"FF803100",
      x"FF863600",
      x"FF8F3E04",
      x"FF914001",
      x"FF954101",
      x"FF944001",
      x"FF933F01",
      x"FF913D01",
      x"FF913D00",
      x"FF953F02",
      x"FF943E01",
      x"FF933F01",
      x"FF974202",
      x"FF974201",
      x"FF9A4601",
      x"FF9B4700",
      x"FF9C4801",
      x"FF994501",
      x"FF9D4901",
      x"FF9D4901",
      x"FF984401",
      x"FF883701",
      x"FF853901",
      x"FF8B3C02",
      x"FF8B3B02",
      x"FF873601",
      x"FF8A3A02",
      x"FF813400",
      x"FF873703",
      x"FF853501",
      x"FF843401",
      x"FF843401",
      x"FF883803",
      x"FF863602",
      x"FF843400",
      x"FF893A02",
      x"FF8A3B03",
      x"FF893A02",
      x"FF823301",
      x"FF7F3201",
      x"FF7F3101",
      x"FF833101",
      x"FF823001",
      x"FF802E01",
      x"FF812F01",
      x"FF823001",
      x"FF843203",
      x"FF812F00",
      x"FF833101",
      x"FF8B3A04",
      x"FF883501",
      x"FF8A3802",
      x"FF883700",
      x"FF873504",
      x"FF873302",
      x"FF8C3A02",
      x"FF8E3A00",
      x"FF923E02",
      x"FF8E3B01",
      x"FF873501",
      x"FF823201",
      x"FF853401",
      x"FF8D3B02",
      x"FF903D01",
      x"FF933F00",
      x"FF944002",
      x"FF923E02",
      x"FF8F3B01",
      x"FF903C00",
      x"FF933D02",
      x"FF913B00",
      x"FF923E01",
      x"FF974102",
      x"FF954000",
      x"FF994401",
      x"FF9B4701",
      x"FF9B4601",
      x"FF984301",
      x"FF9D4901",
      x"FF9D4902",
      x"FF984401",
      x"FF883702",
      x"FF853801",
      x"FF8B3C02",
      x"FF8B3A03",
      x"FF873501",
      x"FF8A3904",
      x"FF833301",
      x"FF873703",
      x"FF823200",
      x"FF853504",
      x"FF833302",
      x"FF853501",
      x"FF863603",
      x"FF853501",
      x"FF893A03",
      x"FF8C3D03",
      x"FF893A02",
      x"FF833402",
      x"FF813402",
      x"FF803001",
      x"FF802E00",
      x"FF812F01",
      x"FF7F2D01",
      x"FF812F01",
      x"FF823001",
      x"FF833102",
      x"FF833102",
      x"FF823001",
      x"FF873601",
      x"FF893602",
      x"FF883501",
      x"FF883700",
      x"FF843202",
      x"FF873303",
      x"FF863300",
      x"FF903B01",
      x"FF8F3B01",
      x"FF913E02",
      x"FF873400",
      x"FF843102",
      x"FF873402",
      x"FF8E3801",
      x"FF903A00",
      x"FF943F01",
      x"FF933D01",
      x"FF923C01",
      x"FF903A01",
      x"FF8F3B01",
      x"FF913B01",
      x"FF903A00",
      x"FF913D01",
      x"FF954001",
      x"FF954000",
      x"FF984300",
      x"FF9A4601",
      x"FF9C4501",
      x"FF9A4301",
      x"FF9D4601",
      x"FF9D4601",
      x"FF974302",
      x"FF853401",
      x"FF833701",
      x"FF8A3B02",
      x"FF893801",
      x"FF873401",
      x"FF893703",
      x"FF833301",
      x"FF863603",
      x"FF823201",
      x"FF853504",
      x"FF823201",
      x"FF843401",
      x"FF843402",
      x"FF863603",
      x"FF843500",
      x"FF893A02",
      x"FF863701",
      x"FF813201",
      x"FF7E3001",
      x"FF823102",
      x"FF7E2D01",
      x"FF823103",
      x"FF7F2E02",
      x"FF7F2E01",
      x"FF802F02",
      x"FF813001",
      x"FF7F2E00",
      x"FF812F02",
      x"FF853302",
      x"FF8C3702",
      x"FF873102",
      x"FF8B3602",
      x"FF843100",
      x"FF843200",
      x"FF853201",
      x"FF8B3701",
      x"FF8C3701",
      x"FF903C03",
      x"FF873501",
      x"FF843002",
      x"FF853101",
      x"FF8D3702",
      x"FF8F3A02",
      x"FF933D02",
      x"FF913B01",
      x"FF923C00",
      x"FF8F3901",
      x"FF8F3802",
      x"FF903901",
      x"FF913B01",
      x"FF923C01",
      x"FF974201",
      x"FF964100",
      x"FF9B4401",
      x"FF9E4704",
      x"FF9D4602",
      x"FF963E00",
      x"FF9D4502",
      x"FF9D4600",
      x"FF964103",
      x"FF843201",
      x"FF853502",
      x"FF8C3C03",
      x"FF8A3803",
      x"FF853401",
      x"FF8A3701",
      x"FF823301",
      x"FF853501",
      x"FF823201",
      x"FF823403",
      x"FF7C2E01",
      x"FF833303",
      x"FF823202",
      x"FF863404",
      x"FF873502",
      x"FF863602",
      x"FF853505",
      x"FF7F2E01",
      x"FF802F01",
      x"FF843302",
      x"FF7E2B01",
      x"FF812F02",
      x"FF812E02",
      x"FF7F2C00",
      x"FF802D01",
      x"FF802E00",
      x"FF802E00",
      x"FF802F01",
      x"FF823001",
      x"FF8E3803",
      x"FF863000",
      x"FF8C3703",
      x"FF853200",
      x"FF863402",
      x"FF853201",
      x"FF8C3602",
      x"FF8B3500",
      x"FF903C02",
      x"FF863401",
      x"FF822E00",
      x"FF833000",
      x"FF8C3701",
      x"FF903B03",
      x"FF933D03",
      x"FF923C01",
      x"FF933D02",
      x"FF913B02",
      x"FF8F3A03",
      x"FF913C02",
      x"FF913D01",
      x"FF923E00",
      x"FF974202",
      x"FF954000",
      x"FF994200",
      x"FF9C4502",
      x"FF9B4400",
      x"FF963E00",
      x"FF9C4403",
      x"FF9A4300",
      x"FF964103",
      x"FF853201",
      x"FF833201",
      x"FF8D3B03",
      x"FF8A3803",
      x"FF853401",
      x"FF893701",
      x"FF823301",
      x"FF873402",
      x"FF823000",
      x"FF853404",
      x"FF802F01",
      x"FF813001",
      x"FF803001",
      x"FF823000",
      x"FF843202",
      x"FF853502",
      x"FF803001",
      x"FF7F2E00",
      x"FF802F00",
      x"FF833202",
      x"FF7F2C02",
      x"FF7F2C00",
      x"FF812E02",
      x"FF7F2C01",
      x"FF812E02",
      x"FF823001",
      x"FF812F01",
      x"FF813000",
      x"FF812D00",
      x"FF8C3602",
      x"FF893302",
      x"FF8C3603",
      x"FF843200",
      x"FF843201",
      x"FF853200",
      x"FF8C3503",
      x"FF8C3501",
      x"FF913B02",
      x"FF8A3701",
      x"FF843001",
      x"FF853101",
      x"FF8C3701",
      x"FF8E3901",
      x"FF923C01",
      x"FF933D01",
      x"FF923C01",
      x"FF8F3901",
      x"FF8E3902",
      x"FF8E3901",
      x"FF903B01",
      x"FF913D01",
      x"FF964102",
      x"FF964101",
      x"FF994101",
      x"FF994201",
      x"FF9C4501",
      x"FF953D00",
      x"FF9B4303",
      x"FF9A4301",
      x"FF954003",
      x"FF843202",
      x"FF833000",
      x"FF8E3903",
      x"FF883502",
      x"FF863402",
      x"FF8A3703",
      x"FF823201",
      x"FF853301",
      x"FF843102",
      x"FF863404",
      x"FF823002",
      x"FF813001",
      x"FF813001",
      x"FF833102",
      x"FF853303",
      x"FF823201",
      x"FF813001",
      x"FF813002",
      x"FF823202",
      x"FF823002",
      x"FF7E2D02",
      x"FF7D2C00",
      x"FF802F02",
      x"FF822E03",
      x"FF802C01",
      x"FF832F01",
      x"FF843002",
      x"FF812F00",
      x"FF812D01",
      x"FF893301",
      x"FF893301",
      x"FF8A3402",
      x"FF883502",
      x"FF843201",
      x"FF873402",
      x"FF8C3404",
      x"FF8C3501",
      x"FF903B01",
      x"FF8D3902",
      x"FF853102",
      x"FF863201",
      x"FF8C3601",
      x"FF8D3801",
      x"FF923C02",
      x"FF943E02",
      x"FF953F03",
      x"FF913B03",
      x"FF8E3703",
      x"FF8D3601",
      x"FF903902",
      x"FF903A01",
      x"FF923D00",
      x"FF943F00",
      x"FF973F01",
      x"FF9A4202",
      x"FF9B4401",
      x"FF943C00",
      x"FF994102",
      x"FF984000",
      x"FF933E02",
      x"FF853203",
      x"FF833100",
      x"FF8C3602",
      x"FF883502",
      x"FF863402",
      x"FF883501",
      x"FF802F00",
      x"FF853301",
      x"FF823001",
      x"FF823101",
      x"FF802F01",
      x"FF7F2E01",
      x"FF7F2E00",
      x"FF833102",
      x"FF833101",
      x"FF823201",
      x"FF802F01",
      x"FF823102",
      x"FF802F00",
      x"FF7F2D02",
      x"FF7F2C02",
      x"FF7C2901",
      x"FF7D2A02",
      x"FF7F2C01",
      x"FF7F2C00",
      x"FF802C01",
      x"FF822E00",
      x"FF822E01",
      x"FF7F2C01",
      x"FF833003",
      x"FF893302",
      x"FF893302",
      x"FF8A3502",
      x"FF833000",
      x"FF873403",
      x"FF8A3401",
      x"FF8B3601",
      x"FF8F3802",
      x"FF913B03",
      x"FF873101",
      x"FF873101",
      x"FF8B3601",
      x"FF8C3701",
      x"FF913C02",
      x"FF933E03",
      x"FF933E02",
      x"FF903B01",
      x"FF8F3A03",
      x"FF8E3701",
      x"FF923901",
      x"FF913600",
      x"FF953C02",
      x"FF953C02",
      x"FF973F01",
      x"FF9A4202",
      x"FF9A4202",
      x"FF953C00",
      x"FF9A4203",
      x"FF994101",
      x"FF923C02",
      x"FF843201",
      x"FF833202",
      x"FF893501",
      x"FF893302",
      x"FF863101",
      x"FF873301",
      x"FF802D01",
      x"FF833100",
      x"FF833100",
      x"FF853304",
      x"FF7F2D01",
      x"FF802F02",
      x"FF813000",
      x"FF823201",
      x"FF813101",
      x"FF7F2E01",
      x"FF813001",
      x"FF802F01",
      x"FF7E2D01",
      x"FF7A2B02",
      x"FF7E2B01",
      x"FF7C2902",
      x"FF7C2901",
      x"FF812E03",
      x"FF802D00",
      x"FF7F2B00",
      x"FF843002",
      x"FF822E01",
      x"FF7F2C02",
      x"FF812E01",
      x"FF8B3503",
      x"FF862F01",
      x"FF8C3603",
      x"FF843001",
      x"FF873403",
      x"FF883200",
      x"FF8C3701",
      x"FF8A3300",
      x"FF903903",
      x"FF873101",
      x"FF863001",
      x"FF8E3803",
      x"FF8C3700",
      x"FF903801",
      x"FF923A02",
      x"FF933B02",
      x"FF903801",
      x"FF8E3501",
      x"FF8E3500",
      x"FF903901",
      x"FF923B02",
      x"FF973F01",
      x"FF943B00",
      x"FF983F02",
      x"FF984001",
      x"FF9B4302",
      x"FF943C00",
      x"FF9A4202",
      x"FF994101",
      x"FF913B02",
      x"FF853302",
      x"FF823002",
      x"FF8A3601",
      x"FF893302",
      x"FF863001",
      x"FF883301",
      x"FF822F01",
      x"FF823001",
      x"FF823000",
      x"FF833002",
      x"FF7E2B01",
      x"FF802F02",
      x"FF813001",
      x"FF813001",
      x"FF7F2E01",
      x"FF7F2E01",
      x"FF823103",
      x"FF813003",
      x"FF7D2C02",
      x"FF7B2C04",
      x"FF7F2C02",
      x"FF7D2A02",
      x"FF7D2A02",
      x"FF802C02",
      x"FF802C00",
      x"FF832D01",
      x"FF832C00",
      x"FF812D01",
      x"FF7F2C01",
      x"FF802D00",
      x"FF8A3402",
      x"FF872F01",
      x"FF8C3503",
      x"FF862F00",
      x"FF873202",
      x"FF863001",
      x"FF8A3401",
      x"FF883000",
      x"FF8D3602",
      x"FF873303",
      x"FF842E00",
      x"FF8A3301",
      x"FF8E3701",
      x"FF913901",
      x"FF933B03",
      x"FF913A01",
      x"FF8F3701",
      x"FF8F3401",
      x"FF8E3401",
      x"FF8F3802",
      x"FF903A03",
      x"FF973F02",
      x"FF983F02",
      x"FF963E01",
      x"FF994101",
      x"FF9A4202",
      x"FF953C00",
      x"FF994102",
      x"FF984001",
      x"FF903801",
      x"FF842F01",
      x"FF802C01",
      x"FF8A3402",
      x"FF883202",
      x"FF893303",
      x"FF873301",
      x"FF822E01",
      x"FF833003",
      x"FF823001",
      x"FF7E2C01",
      x"FF7F2C04",
      x"FF802D01",
      x"FF812F01",
      x"FF812F01",
      x"FF7F2C01",
      x"FF7E2D02",
      x"FF7E2D01",
      x"FF7E2D01",
      x"FF7B2901",
      x"FF782601",
      x"FF7D2A01",
      x"FF7E2B03",
      x"FF7B2801",
      x"FF7B2700",
      x"FF863203",
      x"FF852E01",
      x"FF842D01",
      x"FF832F02",
      x"FF7F2C01",
      x"FF7F2C00",
      x"FF893302",
      x"FF893101",
      x"FF8A3201",
      x"FF862F01",
      x"FF883202",
      x"FF863002",
      x"FF883201",
      x"FF8A3202",
      x"FF8C3402",
      x"FF853102",
      x"FF822C01",
      x"FF8A3302",
      x"FF8F3601",
      x"FF8F3A00",
      x"FF913C01",
      x"FF923D01",
      x"FF8E3900",
      x"FF8E3501",
      x"FF8D3401",
      x"FF8F3601",
      x"FF8E3701",
      x"FF943B02",
      x"FF943B01",
      x"FF963E01",
      x"FF994101",
      x"FF983F01",
      x"FF933A00",
      x"FF973E03",
      x"FF963E01",
      x"FF913802",
      x"FF842F01",
      x"FF822D02",
      x"FF8C3503",
      x"FF883202",
      x"FF873101",
      x"FF883301",
      x"FF843002",
      x"FF7F2C01",
      x"FF812F02",
      x"FF7C2901",
      x"FF7D2A03",
      x"FF812E02",
      x"FF823001",
      x"FF802D01",
      x"FF7D2A01",
      x"FF7D2B01",
      x"FF7E2D01",
      x"FF7C2B00",
      x"FF7B2901",
      x"FF792701",
      x"FF7B2A01",
      x"FF7B2902",
      x"FF7A2802",
      x"FF782401",
      x"FF822F02",
      x"FF873301",
      x"FF832C01",
      x"FF822E00",
      x"FF812D02",
      x"FF822C01",
      x"FF872F02",
      x"FF893202",
      x"FF893001",
      x"FF8A3100",
      x"FF852E01",
      x"FF893102",
      x"FF883001",
      x"FF893101",
      x"FF8A3202",
      x"FF893203",
      x"FF852C00",
      x"FF8B3302",
      x"FF903602",
      x"FF903902",
      x"FF913B01",
      x"FF933D02",
      x"FF8E3701",
      x"FF903B02",
      x"FF8D3701",
      x"FF903602",
      x"FF8F3500",
      x"FF963D01",
      x"FF943C00",
      x"FF953C01",
      x"FF984000",
      x"FF994101",
      x"FF943C00",
      x"FF953A01",
      x"FF973D00",
      x"FF8F3702",
      x"FF862F01",
      x"FF832D00",
      x"FF8B3502",
      x"FF883003",
      x"FF863001",
      x"FF893304",
      x"FF822E01",
      x"FF7F2C00",
      x"FF843002",
      x"FF7B2801",
      x"FF7E2D02",
      x"FF852E01",
      x"FF822E00",
      x"FF7F2D01",
      x"FF7B2902",
      x"FF7B2901",
      x"FF7C2A02",
      x"FF7A2800",
      x"FF7A2800",
      x"FF772401",
      x"FF7D2A01",
      x"FF7B2701",
      x"FF7A2601",
      x"FF7A2602",
      x"FF7D2A00",
      x"FF893404",
      x"FF842D01",
      x"FF832D01",
      x"FF802C01",
      x"FF802B01",
      x"FF852E02",
      x"FF883102",
      x"FF882F01",
      x"FF8C3302",
      x"FF842D01",
      x"FF893103",
      x"FF852D00",
      x"FF8B3303",
      x"FF872F02",
      x"FF893303",
      x"FF852C00",
      x"FF8A3201",
      x"FF8E3401",
      x"FF903602",
      x"FF933A01",
      x"FF943B03",
      x"FF913702",
      x"FF8F3601",
      x"FF8D3401",
      x"FF8F3503",
      x"FF8F3501",
      x"FF953C01",
      x"FF963D01",
      x"FF953C01",
      x"FF994102",
      x"FF984001",
      x"FF953C01",
      x"FF943901",
      x"FF973D02",
      x"FF8E3601",
      x"FF852E00",
      x"FF842E00",
      x"FF8B3602",
      x"FF862E01",
      x"FF852F01",
      x"FF883203",
      x"FF832F01",
      x"FF812D01",
      x"FF822E00",
      x"FF7C2A01",
      x"FF822F03",
      x"FF852F01",
      x"FF822E01",
      x"FF7C2900",
      x"FF792701",
      x"FF7B2903",
      x"FF7C2A04",
      x"FF7B2903",
      x"FF792701",
      x"FF762902",
      x"FF7B2701",
      x"FF792500",
      x"FF782401",
      x"FF792500",
      x"FF7B2701",
      x"FF842F02",
      x"FF862F02",
      x"FF832C01",
      x"FF802A01",
      x"FF802B01",
      x"FF832C01",
      x"FF873001",
      x"FF892F01",
      x"FF8D3402",
      x"FF852E01",
      x"FF872F02",
      x"FF862E01",
      x"FF893102",
      x"FF893102",
      x"FF893302",
      x"FF852C00",
      x"FF883000",
      x"FF8D3301",
      x"FF903602",
      x"FF923801",
      x"FF923901",
      x"FF8F3501",
      x"FF8E3301",
      x"FF8D3201",
      x"FF8D3301",
      x"FF8F3501",
      x"FF923901",
      x"FF943C00",
      x"FF943B01",
      x"FF963E01",
      x"FF963C00",
      x"FF943A01",
      x"FF933A02",
      x"FF973E03",
      x"FF8D3401",
      x"FF822A00",
      x"FF832C01",
      x"FF893302",
      x"FF862D01",
      x"FF842D00",
      x"FF852E01",
      x"FF822E01",
      x"FF802901",
      x"FF822D01",
      x"FF7B2900",
      x"FF812C01",
      x"FF863001",
      x"FF802C01",
      x"FF7A2701",
      x"FF782601",
      x"FF792702",
      x"FF792701",
      x"FF782600",
      x"FF772600",
      x"FF762A01",
      x"FF7D2802",
      x"FF7B2502",
      x"FF792300",
      x"FF7A2601",
      x"FF7C2702",
      x"FF812B02",
      x"FF852F01",
      x"FF842C02",
      x"FF802A01",
      x"FF802B02",
      x"FF802C00",
      x"FF872F01",
      x"FF8A3002",
      x"FF8B3202",
      x"FF852D01",
      x"FF842B01",
      x"FF852D01",
      x"FF883001",
      x"FF893102",
      x"FF893301",
      x"FF852C00",
      x"FF883001",
      x"FF903603",
      x"FF903401",
      x"FF943903",
      x"FF933802",
      x"FF903401",
      x"FF903301",
      x"FF8E3201",
      x"FF903602",
      x"FF903601",
      x"FF913801",
      x"FF953D00",
      x"FF943B01",
      x"FF963D02",
      x"FF973D01",
      x"FF943901",
      x"FF923902",
      x"FF943B01",
      x"FF8A3102",
      x"FF812801",
      x"FF812902",
      x"FF883103",
      x"FF862D02",
      x"FF832C01",
      x"FF852E02",
      x"FF822E01",
      x"FF7F2602",
      x"FF802B02",
      x"FF7B2901",
      x"FF822B02",
      x"FF863001",
      x"FF802C01",
      x"FF7A2602",
      x"FF782601",
      x"FF792702",
      x"FF782601",
      x"FF792702",
      x"FF792701",
      x"FF7A2801",
      x"FF7D2801",
      x"FF7E2902",
      x"FF7E2900",
      x"FF7B2702",
      x"FF7B2800",
      x"FF7F2B01",
      x"FF873303",
      x"FF852D00",
      x"FF802B00",
      x"FF802B02",
      x"FF7F2A02",
      x"FF832B02",
      x"FF872E03",
      x"FF872E01",
      x"FF892F01",
      x"FF842B00",
      x"FF892F03",
      x"FF892E02",
      x"FF892D01",
      x"FF8C3103",
      x"FF882D00",
      x"FF8C3103",
      x"FF903602",
      x"FF8F3401",
      x"FF933802",
      x"FF943903",
      x"FF903501",
      x"FF903401",
      x"FF903402",
      x"FF8E3201",
      x"FF903500",
      x"FF923701",
      x"FF963C01",
      x"FF933801",
      x"FF943A00",
      x"FF973A01",
      x"FF953A03",
      x"FF953A02",
      x"FF953D01",
      x"FF893202",
      x"FF7F2B01",
      x"FF812C01",
      x"FF893303",
      x"FF852D01",
      x"FF862D01",
      x"FF842F01",
      x"FF822E03",
      x"FF7F2901",
      x"FF7D2A00",
      x"FF7D2901",
      x"FF852E01",
      x"FF832E00",
      x"FF7F2B02",
      x"FF7A2601",
      x"FF792500",
      x"FF7B2702",
      x"FF792601",
      x"FF782502",
      x"FF772401",
      x"FF7B2702",
      x"FF7E2902",
      x"FF7E2902",
      x"FF7D2800",
      x"FF7C2802",
      x"FF7C2801",
      x"FF7E2902",
      x"FF863203",
      x"FF852D00",
      x"FF802B01",
      x"FF7F2A01",
      x"FF7E2902",
      x"FF812901",
      x"FF852D01",
      x"FF852C00",
      x"FF8A3102",
      x"FF832D01",
      x"FF862F02",
      x"FF852D02",
      x"FF862D01",
      x"FF8C3103",
      x"FF8B3001",
      x"FF8A2F01",
      x"FF8D3300",
      x"FF8F3400",
      x"FF923701",
      x"FF923702",
      x"FF903401",
      x"FF8F3302",
      x"FF903402",
      x"FF8C3001",
      x"FF8E3200",
      x"FF903400",
      x"FF953B01",
      x"FF923703",
      x"FF923701",
      x"FF973A01",
      x"FF943902",
      x"FF933801",
      x"FF953C02",
      x"FF862F01",
      x"FF7E2901",
      x"FF802B01",
      x"FF863001",
      x"FF832D01",
      x"FF842C01",
      x"FF862E02",
      x"FF822B02",
      x"FF822D01",
      x"FF7E2B01",
      x"FF7D2902",
      x"FF852E03",
      x"FF812D00",
      x"FF7E2901",
      x"FF7B2802",
      x"FF7B2701",
      x"FF7F2B03",
      x"FF7A2700",
      x"FF7A2801",
      x"FF792701",
      x"FF7D2903",
      x"FF7C2701",
      x"FF7E2902",
      x"FF7E2901",
      x"FF7D2801",
      x"FF7C2700",
      x"FF7F2702",
      x"FF842E01",
      x"FF852D01",
      x"FF822C02",
      x"FF7E2900",
      x"FF7E2902",
      x"FF802901",
      x"FF842D01",
      x"FF852E01",
      x"FF893202",
      x"FF822E00",
      x"FF822D01",
      x"FF822B00",
      x"FF862E02",
      x"FF8D3204",
      x"FF8C3101",
      x"FF8B3002",
      x"FF8F3501",
      x"FF8F3401",
      x"FF923701",
      x"FF933802",
      x"FF923602",
      x"FF8F3302",
      x"FF8E3201",
      x"FF8C3001",
      x"FF8F3301",
      x"FF8E3301",
      x"FF973C03",
      x"FF903401",
      x"FF923701",
      x"FF983B02",
      x"FF933802",
      x"FF933801",
      x"FF943B03",
      x"FF872F02",
      x"FF822B02",
      x"FF812A02",
      x"FF872F03",
      x"FF832E01",
      x"FF842C01",
      x"FF872F02",
      x"FF822B02",
      x"FF812E00",
      x"FF7E2A00",
      x"FF7B2600",
      x"FF822B01",
      x"FF812D02",
      x"FF7E2902",
      x"FF7A2700",
      x"FF7C2901",
      x"FF822E02",
      x"FF7E2A00",
      x"FF7B2801",
      x"FF7B2702",
      x"FF7B2902",
      x"FF7C2701",
      x"FF7C2701",
      x"FF7F2A01",
      x"FF7F2A02",
      x"FF7E2901",
      x"FF822A05",
      x"FF832C01",
      x"FF852D01",
      x"FF832E03",
      x"FF7E2900",
      x"FF7E2902",
      x"FF7F2A01",
      x"FF812B00",
      x"FF863002",
      x"FF883101",
      x"FF842D00",
      x"FF832C01",
      x"FF852D01",
      x"FF872F02",
      x"FF8A2F02",
      x"FF8B3101",
      x"FF8A2F01",
      x"FF8D3300",
      x"FF903501",
      x"FF923702",
      x"FF913600",
      x"FF913602",
      x"FF8E3200",
      x"FF8F3301",
      x"FF8E3201",
      x"FF8F3300",
      x"FF903401",
      x"FF963B02",
      x"FF913501",
      x"FF923701",
      x"FF983B02",
      x"FF933802",
      x"FF923702",
      x"FF933A04",
      x"FF862E01",
      x"FF812902",
      x"FF802801",
      x"FF882F03",
      x"FF862D01",
      x"FF842B01",
      x"FF832E00",
      x"FF7E2B01",
      x"FF7F2C01",
      x"FF7D2800",
      x"FF812A03",
      x"FF832F01",
      x"FF812D02",
      x"FF7D2801",
      x"FF7A2700",
      x"FF7E2B01",
      x"FF822E01",
      x"FF7F2A01",
      x"FF7C2801",
      x"FF792501",
      x"FF772500",
      x"FF7E2903",
      x"FF7E2901",
      x"FF7F2B00",
      x"FF802D02",
      x"FF7E2902",
      x"FF802C00",
      x"FF832C01",
      x"FF862E01",
      x"FF852F01",
      x"FF7F2900",
      x"FF7D2804",
      x"FF832A03",
      x"FF842B02",
      x"FF852D01",
      x"FF863101",
      x"FF872D02",
      x"FF872C01",
      x"FF882D02",
      x"FF8A2F01",
      x"FF892E01",
      x"FF8C3102",
      x"FF8B3003",
      x"FF8C3103",
      x"FF903501",
      x"FF913601",
      x"FF913602",
      x"FF913502",
      x"FF8E3201",
      x"FF8E3202",
      x"FF8E3201",
      x"FF8E3201",
      x"FF8E3301",
      x"FF953802",
      x"FF933601",
      x"FF943A01",
      x"FF973D01",
      x"FF953A02",
      x"FF933702",
      x"FF943902",
      x"FF892E02",
      x"FF7D2802",
      x"FF7E2601",
      x"FF893003",
      x"FF832901",
      x"FF852B01",
      x"FF7E2901",
      x"FF7E2A00",
      x"FF822B03",
      x"FF7B2601",
      x"FF7F2A02",
      x"FF822B01",
      x"FF822A01",
      x"FF7E2903",
      x"FF7B2801",
      x"FF802E02",
      x"FF833001",
      x"FF812D02",
      x"FF792402",
      x"FF752101",
      x"FF792600",
      x"FF7F2B02",
      x"FF802B01",
      x"FF7E2901",
      x"FF7E2B01",
      x"FF7C2701",
      x"FF7F2B01",
      x"FF812A00",
      x"FF883003",
      x"FF862E02",
      x"FF822A01",
      x"FF7F2803",
      x"FF802702",
      x"FF832801",
      x"FF872B01",
      x"FF882E01",
      x"FF8A2F02",
      x"FF872C01",
      x"FF892E02",
      x"FF892E01",
      x"FF8A2F02",
      x"FF8C3102",
      x"FF8A2F02",
      x"FF8C3103",
      x"FF903402",
      x"FF903401",
      x"FF913502",
      x"FF913502",
      x"FF8E3201",
      x"FF8E3202",
      x"FF8D3100",
      x"FF8D3100",
      x"FF8F3401",
      x"FF963903",
      x"FF933601",
      x"FF953B03",
      x"FF963C00",
      x"FF943901",
      x"FF923601",
      x"FF933802",
      x"FF882E01",
      x"FF7F2903",
      x"FF802801",
      x"FF872E03",
      x"FF842B00",
      x"FF862D02",
      x"FF7D2800",
      x"FF7E2901",
      x"FF832C04",
      x"FF792401",
      x"FF7F2A02",
      x"FF822B01",
      x"FF802901",
      x"FF7C2702",
      x"FF7A2701",
      x"FF7F2C01",
      x"FF842E02",
      x"FF822A00",
      x"FF7E2703",
      x"FF7B2702",
      x"FF7D2A04",
      x"FF7E2901",
      x"FF7F2B01",
      x"FF7F2A02",
      x"FF7C2900",
      x"FF7C2701",
      x"FF802B01",
      x"FF822A01",
      x"FF882E03",
      x"FF842B00",
      x"FF842C02",
      x"FF7F2702",
      x"FF802802",
      x"FF832801",
      x"FF862A01",
      x"FF872C01",
      x"FF8A2F01",
      x"FF872C00",
      x"FF892E02",
      x"FF892E01",
      x"FF882D01",
      x"FF8B3002",
      x"FF892E01",
      x"FF8B3001",
      x"FF903402",
      x"FF913502",
      x"FF903401",
      x"FF903401",
      x"FF8F3304",
      x"FF8D3102",
      x"FF8C3001",
      x"FF8E3203",
      x"FF8D3301",
      x"FF953903",
      x"FF933600",
      x"FF933901",
      x"FF943A00",
      x"FF923601",
      x"FF8F3401",
      x"FF943904",
      x"FF882E01",
      x"FF7D2701",
      x"FF812802",
      x"FF832A02",
      x"FF832B00",
      x"FF862E03",
      x"FF7C2600",
      x"FF7F2701",
      x"FF812901",
      x"FF7A2501",
      x"FF802B03",
      x"FF812A01",
      x"FF7B2500",
      x"FF792502",
      x"FF7A2700",
      x"FF802C01",
      x"FF832A00",
      x"FF872E03",
      x"FF7E2803",
      x"FF7B2802",
      x"FF7C2903",
      x"FF7E2902",
      x"FF7F2A03",
      x"FF812D02",
      x"FF7D2A02",
      x"FF7C2702",
      x"FF7F2A02",
      x"FF812901",
      x"FF872C02",
      x"FF852C01",
      x"FF862D03",
      x"FF802701",
      x"FF7F2A02",
      x"FF822901",
      x"FF862C01",
      x"FF882E01",
      x"FF8A2F00",
      x"FF872C00",
      x"FF872C01",
      x"FF882D02",
      x"FF892E01",
      x"FF8C3103",
      x"FF872C00",
      x"FF8A2F02",
      x"FF903403",
      x"FF8F3302",
      x"FF8E3201",
      x"FF8D3101",
      x"FF8D3102",
      x"FF8C3001",
      x"FF8B2F00",
      x"FF8C3001",
      x"FF8D3201",
      x"FF943802",
      x"FF933600",
      x"FF933901",
      x"FF943A00",
      x"FF923601",
      x"FF8E3300",
      x"FF913602",
      x"FF872D01",
      x"FF7F2901",
      x"FF812802",
      x"FF812703",
      x"FF812901",
      x"FF842C02",
      x"FF7F2800",
      x"FF832B02",
      x"FF812901",
      x"FF7B2602",
      x"FF7F2A02",
      x"FF812A01",
      x"FF7D2803",
      x"FF782401",
      x"FF7B2701",
      x"FF822D02",
      x"FF873103",
      x"FF802A01",
      x"FF772200",
      x"FF742301",
      x"FF792701",
      x"FF7C2701",
      x"FF802A04",
      x"FF842B01",
      x"FF822902",
      x"FF7D2702",
      x"FF7E2902",
      x"FF852C02",
      x"FF832A02",
      x"FF872E03",
      x"FF852C00",
      x"FF812601",
      x"FF7F2601",
      x"FF832A01",
      x"FF872D01",
      x"FF872C00",
      x"FF8A2F01",
      x"FF872B01",
      x"FF892E01",
      x"FF882D01",
      x"FF893102",
      x"FF8C3102",
      x"FF872C00",
      x"FF8A2D01",
      x"FF8D3101",
      x"FF8E3200",
      x"FF8E3201",
      x"FF8E3202",
      x"FF8C3002",
      x"FF8B2E02",
      x"FF8B2E02",
      x"FF8D3102",
      x"FF8F3000",
      x"FF953702",
      x"FF933501",
      x"FF953701",
      x"FF983B01",
      x"FF953701",
      x"FF8F3300",
      x"FF913502",
      x"FF852B02",
      x"FF7F2902",
      x"FF822A01",
      x"FF822901",
      x"FF7E2502",
      x"FF852C04",
      x"FF812702",
      x"FF832A02",
      x"FF7E2901",
      x"FF7E2901",
      x"FF802B02",
      x"FF7F2B00",
      x"FF7D2801",
      x"FF782401",
      x"FF7B2601",
      x"FF822B00",
      x"FF862E02",
      x"FF782500",
      x"FF762201",
      x"FF752400",
      x"FF752400",
      x"FF7C2701",
      x"FF7D2701",
      x"FF842C03",
      x"FF832A02",
      x"FF7C2601",
      x"FF7C2701",
      x"FF842B02",
      x"FF7F2700",
      x"FF852D03",
      x"FF852C01",
      x"FF842A02",
      x"FF7F2701",
      x"FF822901",
      x"FF852C01",
      x"FF862C00",
      x"FF8B3102",
      x"FF872C02",
      x"FF882D01",
      x"FF892E02",
      x"FF893102",
      x"FF8B3002",
      x"FF872C00",
      x"FF8A2D01",
      x"FF8D3101",
      x"FF8E3200",
      x"FF8F3301",
      x"FF8F3303",
      x"FF8C3001",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8C3001",
      x"FF8D3100",
      x"FF933802",
      x"FF923702",
      x"FF943902",
      x"FF973A00",
      x"FF953702",
      x"FF903501",
      x"FF8F3402",
      x"FF852B02",
      x"FF802802",
      x"FF842901",
      x"FF842A03",
      x"FF802602",
      x"FF832A02",
      x"FF7F2501",
      x"FF832A01",
      x"FF822A04",
      x"FF822A03",
      x"FF812901",
      x"FF822A01",
      x"FF7E2902",
      x"FF782400",
      x"FF7C2702",
      x"FF832C01",
      x"FF832D01",
      x"FF7E2B01",
      x"FF7F2903",
      x"FF7C2601",
      x"FF7A2501",
      x"FF7F2901",
      x"FF7C2700",
      x"FF822A02",
      x"FF812900",
      x"FF7D2701",
      x"FF7B2600",
      x"FF832902",
      x"FF802903",
      x"FF822B02",
      x"FF842C00",
      x"FF832A02",
      x"FF7F2701",
      x"FF802800",
      x"FF842C03",
      x"FF842B01",
      x"FF893101",
      x"FF872C02",
      x"FF872C01",
      x"FF8B2E03",
      x"FF882F01",
      x"FF8B3002",
      x"FF882D01",
      x"FF8A2D01",
      x"FF8D3101",
      x"FF8F3301",
      x"FF903402",
      x"FF8F3303",
      x"FF8E3203",
      x"FF8B2E02",
      x"FF8A2D01",
      x"FF8C3002",
      x"FF8C3000",
      x"FF903500",
      x"FF923702",
      x"FF943902",
      x"FF973C01",
      x"FF923701",
      x"FF8E3300",
      x"FF903603",
      x"FF842B02",
      x"FF7D2902",
      x"FF802900",
      x"FF802801",
      x"FF7E2401",
      x"FF852C04",
      x"FF802601",
      x"FF822901",
      x"FF7C2400",
      x"FF802802",
      x"FF812903",
      x"FF802801",
      x"FF7C2701",
      x"FF782400",
      x"FF7E2903",
      x"FF863002",
      x"FF822B00",
      x"FF822D01",
      x"FF842B02",
      x"FF812B02",
      x"FF7E2602",
      x"FF812B02",
      x"FF7F2901",
      x"FF7E2900",
      x"FF842C01",
      x"FF7E2802",
      x"FF7B2601",
      x"FF812801",
      x"FF7E2803",
      x"FF7F2800",
      x"FF842D01",
      x"FF842C03",
      x"FF7E2802",
      x"FF7E2700",
      x"FF812902",
      x"FF812801",
      x"FF883001",
      x"FF862B02",
      x"FF882C01",
      x"FF882B02",
      x"FF883001",
      x"FF8D3204",
      x"FF872C00",
      x"FF892C01",
      x"FF8E3202",
      x"FF8E3200",
      x"FF8F3301",
      x"FF8D3101",
      x"FF8D3102",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8C3002",
      x"FF8D3201",
      x"FF903701",
      x"FF913702",
      x"FF923901",
      x"FF953B01",
      x"FF913600",
      x"FF8D3300",
      x"FF8E3401",
      x"FF822800",
      x"FF7D2600",
      x"FF822901",
      x"FF832902",
      x"FF812703",
      x"FF822902",
      x"FF7F2501",
      x"FF812800",
      x"FF7F2502",
      x"FF802601",
      x"FF812702",
      x"FF812702",
      x"FF7C2602",
      x"FF782401",
      x"FF7E2A02",
      x"FF842D00",
      x"FF812801",
      x"FF842C01",
      x"FF852A00",
      x"FF802A01",
      x"FF7D2702",
      x"FF852C02",
      x"FF812800",
      x"FF7F2602",
      x"FF842C03",
      x"FF7F2702",
      x"FF7B2300",
      x"FF7F2801",
      x"FF7D2902",
      x"FF812701",
      x"FF842D02",
      x"FF873101",
      x"FF842B02",
      x"FF7F2700",
      x"FF832C02",
      x"FF842B01",
      x"FF842D03",
      x"FF822900",
      x"FF852C01",
      x"FF892E03",
      x"FF8A2F01",
      x"FF8D3203",
      x"FF872C00",
      x"FF882D00",
      x"FF8C3002",
      x"FF8D3101",
      x"FF8F3302",
      x"FF8D3102",
      x"FF8C3102",
      x"FF8A2F03",
      x"FF892C01",
      x"FF8B2E02",
      x"FF8D3101",
      x"FF8F3301",
      x"FF923702",
      x"FF923702",
      x"FF943901",
      x"FF923602",
      x"FF8E3201",
      x"FF903403",
      x"FF822801",
      x"FF7D2301",
      x"FF802601",
      x"FF822901",
      x"FF802601",
      x"FF802801",
      x"FF7D2501",
      x"FF7F2502",
      x"FF7F2601",
      x"FF842901",
      x"FF822801",
      x"FF7F2603",
      x"FF7B2601",
      x"FF792400",
      x"FF7F2802",
      x"FF832B03",
      x"FF7F2802",
      x"FF842D01",
      x"FF832B00",
      x"FF832903",
      x"FF7F2703",
      x"FF822900",
      x"FF822902",
      x"FF802602",
      x"FF812901",
      x"FF812903",
      x"FF7C2401",
      x"FF7F2801",
      x"FF7E2902",
      x"FF822902",
      x"FF852E02",
      x"FF893203",
      x"FF842A00",
      x"FF812901",
      x"FF822A02",
      x"FF852C01",
      x"FF862F03",
      x"FF852C02",
      x"FF842B00",
      x"FF882D01",
      x"FF8A2F01",
      x"FF8B3001",
      x"FF872C01",
      x"FF882D00",
      x"FF8C3001",
      x"FF8E3201",
      x"FF8D3100",
      x"FF8C3001",
      x"FF8C3102",
      x"FF8A2F02",
      x"FF882B01",
      x"FF8B2E03",
      x"FF8D3101",
      x"FF903402",
      x"FF923702",
      x"FF913601",
      x"FF943901",
      x"FF913602",
      x"FF8D3100",
      x"FF8F3302",
      x"FF812700",
      x"FF7E2402",
      x"FF7F2501",
      x"FF822901",
      x"FF812802",
      x"FF802901",
      x"FF7F2702",
      x"FF822803",
      x"FF802700",
      x"FF842900",
      x"FF852A02",
      x"FF7E2501",
      x"FF7B2601",
      x"FF7C2600",
      x"FF802801",
      x"FF802801",
      x"FF842B02",
      x"FF862F01",
      x"FF832F01",
      x"FF802B01",
      x"FF7D2601",
      x"FF802700",
      x"FF822803",
      x"FF812702",
      x"FF7F2701",
      x"FF822A03",
      x"FF7A2200",
      x"FF7F2702",
      x"FF7F2801",
      x"FF812901",
      x"FF7F2A00",
      x"FF8B3104",
      x"FF872C00",
      x"FF812801",
      x"FF812801",
      x"FF862B01",
      x"FF832C01",
      x"FF842B02",
      x"FF842B01",
      x"FF8B3002",
      x"FF8A2F00",
      x"FF892F00",
      x"FF882D02",
      x"FF892E01",
      x"FF8B2F01",
      x"FF8D3101",
      x"FF8D3100",
      x"FF8B2F00",
      x"FF8B3001",
      x"FF892E01",
      x"FF892C01",
      x"FF8A2D01",
      x"FF8C3001",
      x"FF8F3301",
      x"FF923702",
      x"FF903500",
      x"FF943901",
      x"FF903401",
      x"FF8B2F00",
      x"FF8E3302",
      x"FF812700",
      x"FF7E2402",
      x"FF802601",
      x"FF812800",
      x"FF822901",
      x"FF822A01",
      x"FF802803",
      x"FF822802",
      x"FF832801",
      x"FF862B01",
      x"FF852C02",
      x"FF7E2802",
      x"FF802803",
      x"FF7F2701",
      x"FF822902",
      x"FF832A00",
      x"FF842B00",
      x"FF872F03",
      x"FF812D01",
      x"FF7F2C02",
      x"FF802A00",
      x"FF812701",
      x"FF822803",
      x"FF802600",
      x"FF7E2600",
      x"FF812901",
      x"FF7E2602",
      x"FF7E2602",
      x"FF822A02",
      x"FF812B02",
      x"FF7E2A01",
      x"FF892F03",
      x"FF8A2F01",
      x"FF842A03",
      x"FF822802",
      x"FF872D02",
      x"FF842E01",
      x"FF852C02",
      x"FF852D02",
      x"FF8F3404",
      x"FF8C3102",
      x"FF8A2F00",
      x"FF872C01",
      x"FF882D01",
      x"FF8C3001",
      x"FF8D3100",
      x"FF8E3201",
      x"FF8C3001",
      x"FF8B3001",
      x"FF892E01",
      x"FF892C01",
      x"FF882B00",
      x"FF8C3000",
      x"FF8F3301",
      x"FF923702",
      x"FF903500",
      x"FF943901",
      x"FF923603",
      x"FF8C3000",
      x"FF8E3202",
      x"FF812701",
      x"FF7E2402",
      x"FF812702",
      x"FF822901",
      x"FF832A01",
      x"FF812A01",
      x"FF802801",
      x"FF812802",
      x"FF832701",
      x"FF862B00",
      x"FF832B01",
      x"FF7D2701",
      x"FF7F2701",
      x"FF7F2700",
      x"FF832A02",
      x"FF832A01",
      x"FF852C01",
      x"FF822901",
      x"FF812902",
      x"FF7F2901",
      x"FF832D01",
      x"FF802A00",
      x"FF7F2901",
      x"FF812903",
      x"FF812801",
      x"FF7D2701",
      x"FF7C2601",
      x"FF7C2603",
      x"FF7F2701",
      x"FF812903",
      x"FF802702",
      x"FF862B01",
      x"FF8A2F01",
      x"FF852C03",
      x"FF812901",
      x"FF852C01",
      x"FF862E01",
      x"FF872E03",
      x"FF862B00",
      x"FF8E3302",
      x"FF8B3001",
      x"FF892E01",
      x"FF872C00",
      x"FF872C00",
      x"FF8B2E02",
      x"FF8D3101",
      x"FF8E3202",
      x"FF8A2E00",
      x"FF8B2E02",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF892C00",
      x"FF8D3101",
      x"FF8F3300",
      x"FF923603",
      x"FF913601",
      x"FF933801",
      x"FF933803",
      x"FF8B3101",
      x"FF8C3202",
      x"FF812703",
      x"FF7D2301",
      x"FF822803",
      x"FF812702",
      x"FF812802",
      x"FF7F2602",
      x"FF7D2701",
      x"FF7E2801",
      x"FF802802",
      x"FF852902",
      x"FF802602",
      x"FF7F2502",
      x"FF802803",
      x"FF822A03",
      x"FF842B03",
      x"FF852C01",
      x"FF862C01",
      x"FF832B01",
      x"FF7F2A02",
      x"FF7C2702",
      x"FF832B01",
      x"FF822D01",
      x"FF7D2801",
      x"FF802802",
      x"FF822A02",
      x"FF7E2700",
      x"FF7C2702",
      x"FF7B2602",
      x"FF822A02",
      x"FF802A01",
      x"FF7F2700",
      x"FF872D03",
      x"FF882E02",
      x"FF822A01",
      x"FF7F2701",
      x"FF832A01",
      x"FF832B02",
      x"FF842B02",
      x"FF842801",
      x"FF892E01",
      x"FF892E01",
      x"FF882D01",
      x"FF882D00",
      x"FF882D01",
      x"FF8A2D01",
      x"FF8C3001",
      x"FF8D3101",
      x"FF8C3001",
      x"FF8B2E02",
      x"FF8A2D01",
      x"FF892C01",
      x"FF8A2D01",
      x"FF8E3202",
      x"FF8E3200",
      x"FF913502",
      x"FF903500",
      x"FF933801",
      x"FF913601",
      x"FF8B3000",
      x"FF8D3202",
      x"FF7F2501",
      x"FF7C2200",
      x"FF802601",
      x"FF7F2500",
      x"FF802601",
      x"FF7F2602",
      x"FF7F2803",
      x"FF7E2901",
      x"FF7F2702",
      x"FF852902",
      x"FF7F2602",
      x"FF7E2502",
      x"FF802802",
      x"FF822902",
      x"FF812801",
      x"FF842A01",
      x"FF852B00",
      x"FF822A01",
      x"FF7D2802",
      x"FF7B2601",
      x"FF802801",
      x"FF812B00",
      x"FF7E2901",
      x"FF7E2600",
      x"FF812900",
      x"FF7F2901",
      x"FF802A04",
      x"FF7B2601",
      x"FF7F2801",
      x"FF802C01",
      x"FF802A01",
      x"FF822901",
      x"FF872E01",
      x"FF812902",
      x"FF7E2702",
      x"FF7F2702",
      x"FF812901",
      x"FF812A00",
      x"FF822901",
      x"FF862C02",
      x"FF872C01",
      x"FF882D02",
      x"FF882D01",
      x"FF882D00",
      x"FF892C01",
      x"FF8C3001",
      x"FF8D3101",
      x"FF8C3001",
      x"FF8C2F03",
      x"FF8B2E02",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8E3201",
      x"FF8E3200",
      x"FF8F3300",
      x"FF8F3400",
      x"FF933801",
      x"FF913500",
      x"FF8A3000",
      x"FF8D3203",
      x"FF812702",
      x"FF7E2401",
      x"FF812703",
      x"FF7F2501",
      x"FF812702",
      x"FF7F2602",
      x"FF7D2702",
      x"FF7E2901",
      x"FF7F2802",
      x"FF842902",
      x"FF7E2601",
      x"FF7D2501",
      x"FF802700",
      x"FF832A02",
      x"FF832801",
      x"FF842801",
      x"FF842A01",
      x"FF822A02",
      x"FF7C2701",
      x"FF7B2602",
      x"FF802702",
      x"FF802A00",
      x"FF7F2A01",
      x"FF7F2701",
      x"FF832B02",
      x"FF812B01",
      x"FF7F2A03",
      x"FF7A2500",
      x"FF7D2802",
      x"FF7D2900",
      x"FF7F2A02",
      x"FF802701",
      x"FF862D01",
      x"FF802A03",
      x"FF7A2501",
      x"FF7C2501",
      x"FF812901",
      x"FF822B01",
      x"FF812801",
      x"FF822901",
      x"FF862A02",
      x"FF872C01",
      x"FF892E02",
      x"FF872C00",
      x"FF892C01",
      x"FF8C3001",
      x"FF8D3101",
      x"FF8C3001",
      x"FF8A2D01",
      x"FF892C00",
      x"FF892C00",
      x"FF8A2E01",
      x"FF8F3302",
      x"FF8F3300",
      x"FF913502",
      x"FF8F3400",
      x"FF933801",
      x"FF933702",
      x"FF8B3101",
      x"FF8D3202",
      x"FF812702",
      x"FF7E2401",
      x"FF822803",
      x"FF7E2401",
      x"FF802701",
      x"FF7E2501",
      x"FF7C2500",
      x"FF7C2700",
      x"FF7E2701",
      x"FF842B02",
      x"FF7C2501",
      x"FF7E2702",
      x"FF832A03",
      x"FF832902",
      x"FF832701",
      x"FF842801",
      x"FF862C02",
      x"FF812802",
      x"FF7A2500",
      x"FF7A2401",
      x"FF7E2501",
      x"FF832C01",
      x"FF812A00",
      x"FF7E2900",
      x"FF822A03",
      x"FF812901",
      x"FF802A01",
      x"FF7B2702",
      x"FF7F2702",
      x"FF7C2700",
      x"FF812C03",
      x"FF822B02",
      x"FF873004",
      x"FF802A01",
      x"FF7A2501",
      x"FF782400",
      x"FF7F2903",
      x"FF812A02",
      x"FF802801",
      x"FF832A01",
      x"FF892E02",
      x"FF872C00",
      x"FF892E01",
      x"FF892E01",
      x"FF892C01",
      x"FF8C3001",
      x"FF8D3100",
      x"FF8C3001",
      x"FF8D3102",
      x"FF8A2E00",
      x"FF8A2D01",
      x"FF8A2E01",
      x"FF903403",
      x"FF903401",
      x"FF913502",
      x"FF913601",
      x"FF943901",
      x"FF923702",
      x"FF8B2F00",
      x"FF8C3003",
      x"FF802701",
      x"FF7A2400",
      x"FF802902",
      x"FF802702",
      x"FF812902",
      x"FF7D2601",
      x"FF7B2602",
      x"FF7A2500",
      x"FF802701",
      x"FF832901",
      x"FF7F2602",
      x"FF812701",
      x"FF842B03",
      x"FF802702",
      x"FF822902",
      x"FF832A02",
      x"FF832B01",
      x"FF7E2902",
      x"FF792400",
      x"FF7A2602",
      x"FF7D2501",
      x"FF832B01",
      x"FF832C00",
      x"FF802901",
      x"FF802801",
      x"FF822A01",
      x"FF802A01",
      x"FF7B2602",
      x"FF7D2501",
      x"FF7F2A03",
      x"FF7E2901",
      x"FF7F2800",
      x"FF862F02",
      x"FF822B02",
      x"FF7C2701",
      x"FF782401",
      x"FF812803",
      x"FF832A02",
      x"FF832A02",
      x"FF842900",
      x"FF882D01",
      x"FF882D01",
      x"FF8A2F02",
      x"FF8B3003",
      x"FF8A2D01",
      x"FF8D3102",
      x"FF8D3100",
      x"FF8C3001",
      x"FF8D3102",
      x"FF8A2E00",
      x"FF882B00",
      x"FF892C00",
      x"FF8F3302",
      x"FF8F3301",
      x"FF913502",
      x"FF913601",
      x"FF923700",
      x"FF923702",
      x"FF8D3100",
      x"FF8A2E01",
      x"FF7F2601",
      x"FF7B2401",
      x"FF7F2802",
      x"FF7F2602",
      x"FF802701",
      x"FF7C2500",
      x"FF7B2501",
      x"FF7A2501",
      x"FF802801",
      x"FF852A02",
      x"FF7F2601",
      x"FF832802",
      x"FF822901",
      x"FF812801",
      x"FF842B03",
      x"FF822902",
      x"FF802800",
      x"FF7B2600",
      x"FF792301",
      x"FF782401",
      x"FF7C2501",
      x"FF862D02",
      x"FF852D00",
      x"FF812901",
      x"FF822A03",
      x"FF822A01",
      x"FF802A01",
      x"FF7A2601",
      x"FF7C2400",
      x"FF802B04",
      x"FF7F2A01",
      x"FF812901",
      x"FF872F02",
      x"FF842C02",
      x"FF7F2902",
      x"FF7A2602",
      x"FF812803",
      x"FF822901",
      x"FF842A02",
      x"FF842900",
      x"FF862B00",
      x"FF872C01",
      x"FF8A2F02",
      x"FF8A2F02",
      x"FF8B2E02",
      x"FF8E3202",
      x"FF8D3101",
      x"FF8D3102",
      x"FF8D3102",
      x"FF8C3001",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8E3201",
      x"FF8E3200",
      x"FF903401",
      x"FF913601",
      x"FF933800",
      x"FF933702",
      x"FF8D3101",
      x"FF8B2F01",
      x"FF802602",
      x"FF7C2402",
      x"FF7E2703",
      x"FF7E2502",
      x"FF802703",
      x"FF7A2300",
      x"FF7A2402",
      x"FF7A2401",
      x"FF822902",
      x"FF842902",
      x"FF7E2501",
      x"FF812601",
      x"FF812801",
      x"FF812801",
      x"FF832A02",
      x"FF822902",
      x"FF822A01",
      x"FF7C2601",
      x"FF782200",
      x"FF762201",
      x"FF7A2300",
      x"FF862C01",
      x"FF842B00",
      x"FF822902",
      x"FF802801",
      x"FF822B01",
      x"FF812B01",
      x"FF7B2702",
      x"FF7C2500",
      x"FF7E2902",
      x"FF7E2901",
      x"FF802901",
      x"FF852D01",
      x"FF842C01",
      x"FF7E2802",
      x"FF7B2601",
      x"FF7E2802",
      x"FF802901",
      x"FF822A02",
      x"FF832A00",
      x"FF872C01",
      x"FF872B01",
      x"FF872C02",
      x"FF862B00",
      x"FF8A2D01",
      x"FF8D3101",
      x"FF8D3101",
      x"FF8B2F01",
      x"FF8C3001",
      x"FF8B2F00",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8E3202",
      x"FF8E3200",
      x"FF913502",
      x"FF923702",
      x"FF933801",
      x"FF933702",
      x"FF8D3101",
      x"FF8B2F02",
      x"FF7E2401",
      x"FF7A2301",
      x"FF7C2601",
      x"FF7D2401",
      x"FF802703",
      x"FF792200",
      x"FF792301",
      x"FF7A2402",
      x"FF822902",
      x"FF832901",
      x"FF7F2602",
      x"FF812601",
      x"FF822901",
      x"FF812801",
      x"FF842B03",
      x"FF822901",
      x"FF812902",
      x"FF7B2502",
      x"FF762000",
      x"FF772301",
      x"FF7E2502",
      x"FF832A02",
      x"FF852D01",
      x"FF822B00",
      x"FF812901",
      x"FF812901",
      x"FF812902",
      x"FF7D2502",
      x"FF792502",
      x"FF7A2501",
      x"FF7D2801",
      x"FF7F2703",
      x"FF832A02",
      x"FF822B02",
      x"FF802803",
      x"FF7C2702",
      x"FF7D2802",
      x"FF7F2802",
      x"FF822901",
      x"FF822901",
      x"FF862A01",
      x"FF862A02",
      x"FF892C02",
      x"FF872A00",
      x"FF892C00",
      x"FF8E3202",
      x"FF8C3001",
      x"FF8C3002",
      x"FF8D3102",
      x"FF8B2F01",
      x"FF8A2D01",
      x"FF892C01",
      x"FF8C3001",
      x"FF8E3201",
      x"FF8F3302",
      x"FF923603",
      x"FF953703",
      x"FF913601",
      x"FF8D3100",
      x"FF882D02",
      x"FF7C2502",
      x"FF7C2401",
      x"FF802804",
      x"FF802601",
      x"FF802703",
      x"FF7A2201",
      x"FF7C2500",
      x"FF7F2703",
      x"FF822B01",
      x"FF802800",
      x"FF802503",
      x"FF812501",
      x"FF7F2601",
      x"FF7F2501",
      x"FF822803",
      x"FF7F2701",
      x"FF7B2600",
      x"FF792202",
      x"FF761F01",
      x"FF792302",
      x"FF7D2401",
      x"FF822C03",
      x"FF842E01",
      x"FF842D01",
      x"FF812A01",
      x"FF812901",
      x"FF812902",
      x"FF7E2603",
      x"FF782401",
      x"FF7B2601",
      x"FF7E2903",
      x"FF7E2602",
      x"FF822901",
      x"FF812A02",
      x"FF7F2702",
      x"FF7D2803",
      x"FF7B2600",
      x"FF802903",
      x"FF822901",
      x"FF822901",
      x"FF852A01",
      x"FF862A02",
      x"FF8A2E02",
      x"FF8A2D02",
      x"FF892C00",
      x"FF8E3202",
      x"FF8C3000",
      x"FF8D3102",
      x"FF8C3001",
      x"FF8B2F01",
      x"FF8B2E02",
      x"FF8A2D01",
      x"FF8C3002",
      x"FF8E3202",
      x"FF8E3201",
      x"FF913503",
      x"FF923401",
      x"FF903500",
      x"FF8D3100",
      x"FF882D02",
      x"FF7C2502",
      x"FF7C2400",
      x"FF7E2602",
      x"FF7F2501",
      x"FF7F2602",
      x"FF7A2301",
      x"FF7E2702",
      x"FF7F2602",
      x"FF832A01",
      x"FF842B02",
      x"FF802603",
      x"FF802701",
      x"FF802802",
      x"FF7F2500",
      x"FF822803",
      x"FF7F2701",
      x"FF7D2802",
      x"FF782201",
      x"FF741D00",
      x"FF782201",
      x"FF7C2400",
      x"FF812C02",
      x"FF862F02",
      x"FF852D02",
      x"FF802901",
      x"FF812901",
      x"FF802801",
      x"FF7D2602",
      x"FF7A2501",
      x"FF7A2400",
      x"FF7C2703",
      x"FF7E2601",
      x"FF822902",
      x"FF832C01",
      x"FF812904",
      x"FF7B2601",
      x"FF7C2701",
      x"FF7E2701",
      x"FF822902",
      x"FF812800",
      x"FF842B00",
      x"FF872D02",
      x"FF892E01",
      x"FF8C3003",
      x"FF8A2D01",
      x"FF8E3202",
      x"FF8C3000",
      x"FF8C3001",
      x"FF8B2F00",
      x"FF892D00",
      x"FF8A2D01",
      x"FF892C00",
      x"FF8D3102",
      x"FF8E3202",
      x"FF8E3201",
      x"FF8F3301",
      x"FF933502",
      x"FF933702",
      x"FF8E3200",
      x"FF882D02",
      x"FF7B2401",
      x"FF7B2300",
      x"FF7E2602",
      x"FF7F2501",
      x"FF802702",
      x"FF7B2301",
      x"FF7C2601",
      x"FF7C2301",
      x"FF852C01",
      x"FF852C01",
      x"FF802602",
      x"FF832A03",
      x"FF812A02",
      x"FF812801",
      x"FF812801",
      x"FF812902",
      x"FF7E2903",
      x"FF792202",
      x"FF772002",
      x"FF792302",
      x"FF7D2601",
      x"FF812901",
      x"FF842A00",
      x"FF872D02",
      x"FF832B02",
      x"FF802801",
      x"FF822A02",
      x"FF7B2301",
      x"FF7B2702",
      x"FF782201",
      x"FF7B2502",
      x"FF7F2701",
      x"FF812801",
      x"FF832C01",
      x"FF812904",
      x"FF7C2702",
      x"FF7C2701",
      x"FF7D2701",
      x"FF812801",
      x"FF802700",
      x"FF842B00",
      x"FF852C00",
      x"FF882E00",
      x"FF8A2F02",
      x"FF892C00",
      x"FF8B2F00",
      x"FF8C3000",
      x"FF8C3001",
      x"FF8B2F00",
      x"FF892D00",
      x"FF8A2D01",
      x"FF892C00",
      x"FF8B2E01",
      x"FF8D3102",
      x"FF8F3302",
      x"FF8F3301",
      x"FF913401",
      x"FF913601",
      x"FF8E3200",
      x"FF882D02",
      x"FF7B2502",
      x"FF7D2502",
      x"FF7E2602",
      x"FF7F2501",
      x"FF7F2602",
      x"FF7A2201",
      x"FF7B2401",
      x"FF812804",
      x"FF882D01",
      x"FF842A01",
      x"FF812802",
      x"FF812A01",
      x"FF802801",
      x"FF832A02",
      x"FF842B03",
      x"FF812902",
      x"FF7E2803",
      x"FF7A2403",
      x"FF782103",
      x"FF782201",
      x"FF7B2500",
      x"FF7E2803",
      x"FF832A01",
      x"FF852C01",
      x"FF842C03",
      x"FF7E2601",
      x"FF822A02",
      x"FF7E2601",
      x"FF7C2702",
      x"FF792400",
      x"FF7F2803",
      x"FF832901",
      x"FF802901",
      x"FF832E01",
      x"FF7F2A00",
      x"FF7F2802",
      x"FF7F2A02",
      x"FF7C2701",
      x"FF7F2802",
      x"FF7F2603",
      x"FF862B01",
      x"FF872C01",
      x"FF882D01",
      x"FF892E02",
      x"FF882D01",
      x"FF8A2F02",
      x"FF8A2F02",
      x"FF8A2F00",
      x"FF8B2E02",
      x"FF892C00",
      x"FF8A2D01",
      x"FF892C01",
      x"FF882D01",
      x"FF8B3002",
      x"FF8D3301",
      x"FF8D3301",
      x"FF8B3202",
      x"FF903503",
      x"FF8D3200",
      x"FF862C02",
      x"FF7D2702",
      x"FF7B2601",
      x"FF7F2701",
      x"FF7E2601",
      x"FF812802",
      x"FF7B2501",
      x"FF7B2501",
      x"FF802701",
      x"FF822901",
      x"FF812801",
      x"FF812801",
      x"FF812800",
      x"FF7F2702",
      x"FF842A00",
      x"FF852900",
      x"FF832A02",
      x"FF7B2402",
      x"FF772200",
      x"FF762101",
      x"FF762101",
      x"FF7D2701",
      x"FF7C2702",
      x"FF842B01",
      x"FF832B01",
      x"FF812901",
      x"FF7F2702",
      x"FF822A02",
      x"FF7F2802",
      x"FF7A2601",
      x"FF782400",
      x"FF7D2702",
      x"FF832A01",
      x"FF822901",
      x"FF842C01",
      x"FF802C01",
      x"FF7C2802",
      x"FF7E2902",
      x"FF7C2600",
      x"FF812902",
      x"FF802803",
      x"FF882C01",
      x"FF882D01",
      x"FF882D01",
      x"FF882D01",
      x"FF882D01",
      x"FF8A2F02",
      x"FF8A2F02",
      x"FF8A2F00",
      x"FF8C2F03",
      x"FF8A2D01",
      x"FF8B2E02",
      x"FF8B2E02",
      x"FF892E02",
      x"FF8C3102",
      x"FF8D3301",
      x"FF8E3402",
      x"FF8B3202",
      x"FF923704",
      x"FF8D3101",
      x"FF842A01",
      x"FF7B2500",
      x"FF7B2601",
      x"FF7C2400",
      x"FF802802",
      x"FF802701",
      x"FF7E2803",
      x"FF7D2702",
      x"FF812903",
      x"FF832A01",
      x"FF832903",
      x"FF812702",
      x"FF812801",
      x"FF7D2500",
      x"FF852B01",
      x"FF862B01",
      x"FF812800",
      x"FF7C2402",
      x"FF772201",
      x"FF752101",
      x"FF772103",
      x"FF7C2501",
      x"FF7D2802",
      x"FF822901",
      x"FF822A01",
      x"FF7F2701",
      x"FF802803",
      x"FF822A01",
      x"FF822A03",
      x"FF7B2702",
      x"FF782401",
      x"FF7D2803",
      x"FF822901",
      x"FF822902",
      x"FF822B01",
      x"FF812D02",
      x"FF7A2601",
      x"FF812903",
      x"FF802801",
      x"FF832A02",
      x"FF822902",
      x"FF872C00",
      x"FF872C01",
      x"FF872C01",
      x"FF882D01",
      x"FF882D01",
      x"FF882D01",
      x"FF8A2F02",
      x"FF892E00",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF882D01",
      x"FF8D3202",
      x"FF8D3300",
      x"FF8F3502",
      x"FF8B3201",
      x"FF913602",
      x"FF8C3001",
      x"FF832901",
      x"FF7C2601",
      x"FF7E2904",
      x"FF7E2600",
      x"FF812903",
      x"FF802702",
      x"FF7D2602",
      x"FF7B2501",
      x"FF812903",
      x"FF842B01",
      x"FF822902",
      x"FF812702",
      x"FF822802",
      x"FF7F2702",
      x"FF852B01",
      x"FF872C01",
      x"FF822901",
      x"FF7C2301",
      x"FF7A2302",
      x"FF772202",
      x"FF772002",
      x"FF7C2300",
      x"FF7C2701",
      x"FF832A01",
      x"FF832B03",
      x"FF802802",
      x"FF7F2701",
      x"FF802800",
      x"FF812A03",
      x"FF7B2802",
      x"FF7A2803",
      x"FF7E2903",
      x"FF812901",
      x"FF7D2700",
      x"FF802B02",
      x"FF812B03",
      x"FF792301",
      x"FF7F2701",
      x"FF802701",
      x"FF872E04",
      x"FF822902",
      x"FF862B01",
      x"FF872C01",
      x"FF872C00",
      x"FF882D01",
      x"FF892E02",
      x"FF872C00",
      x"FF892E01",
      x"FF8A2F00",
      x"FF8B2E02",
      x"FF8B2E02",
      x"FF8A2D01",
      x"FF8A2D01",
      x"FF8A2F02",
      x"FF8D3301",
      x"FF8C3200",
      x"FF8E3400",
      x"FF8C3301",
      x"FF903501",
      x"FF8B2F00",
      x"FF822801",
      x"FF7A2501",
      x"FF7C2702",
      x"FF7D2500",
      x"FF802802",
      x"FF7F2601",
      x"FF7E2803",
      x"FF7B2501",
      x"FF802802",
      x"FF852C02",
      x"FF812801",
      x"FF812702",
      x"FF802601",
      x"FF812903",
      x"FF852B01",
      x"FF862B01",
      x"FF822801",
      x"FF7F2503",
      x"FF782100",
      x"FF772002",
      x"FF771F01",
      x"FF802701",
      x"FF7D2802",
      x"FF802C01",
      x"FF802901",
      x"FF7E2902",
      x"FF7E2901",
      x"FF7D2802",
      x"FF7E2904",
      x"FF7D2803",
      x"FF7D2803",
      x"FF7F2701",
      x"FF822A01",
      x"FF7E2901",
      x"FF812D03",
      x"FF7F2C02",
      x"FF782401",
      x"FF812903",
      x"FF7F2702",
      x"FF872E03",
      x"FF822902",
      x"FF862B01",
      x"FF842800",
      x"FF882C02",
      x"FF872C01",
      x"FF882D01",
      x"FF862B00",
      x"FF892E01",
      x"FF8B3001",
      x"FF8A2F02",
      x"FF892E01",
      x"FF892E01",
      x"FF892E01",
      x"FF8A2F02",
      x"FF8D3203",
      x"FF8F3503",
      x"FF8E3400",
      x"FF8D3301",
      x"FF8F3301",
      x"FF8A2F01",
      x"FF812802",
      x"FF792400",
      x"FF7D2803",
      x"FF7C2400",
      x"FF802602",
      x"FF7E2602",
      x"FF7C2700",
      x"FF7D2801",
      x"FF812902",
      x"FF832902",
      x"FF802500",
      x"FF812900",
      x"FF7E2802",
      x"FF822A02",
      x"FF832A00",
      x"FF832A01",
      x"FF7D2401",
      x"FF7A2400",
      x"FF752001",
      x"FF752002",
      x"FF792302",
      x"FF842901",
      x"FF7C2702",
      x"FF802D01",
      x"FF822B03",
      x"FF7C2701",
      x"FF7E2901",
      x"FF7D2801",
      x"FF7D2802",
      x"FF7D2803",
      x"FF7D2803",
      x"FF802801",
      x"FF852D04",
      x"FF7E2601",
      x"FF822C03",
      x"FF802A01",
      x"FF7C2502",
      x"FF802802",
      x"FF7B2300",
      x"FF883003",
      x"FF842B02",
      x"FF872C02",
      x"FF852A01",
      x"FF862A00",
      x"FF872B01",
      x"FF8A2F03",
      x"FF882D00",
      x"FF892E01",
      x"FF8A2F00",
      x"FF8A2F02",
      x"FF892E01",
      x"FF8A2F02",
      x"FF892E01",
      x"FF8A2F02",
      x"FF8D3203",
      x"FF8D3301",
      x"FF8E3401",
      x"FF8D3301",
      x"FF8F3301",
      x"FF892E00",
      x"FF802702",
      x"FF792400",
      x"FF7B2602",
      x"FF7D2501",
      x"FF812803",
      x"FF7E2602",
      x"FF7C2700",
      x"FF7C2701",
      x"FF812901",
      x"FF7F2801",
      x"FF812701",
      x"FF832A01",
      x"FF7E2501",
      x"FF812901",
      x"FF842B01",
      x"FF842B02",
      x"FF7E2501",
      x"FF792300",
      x"FF762101",
      x"FF752101",
      x"FF792401",
      x"FF822900",
      x"FF7B2701",
      x"FF7E2B01",
      x"FF812B02",
      x"FF7D2802",
      x"FF7F2A02",
      x"FF7F2A01",
      x"FF7C2701",
      x"FF7C2702",
      x"FF7B2601",
      x"FF802801",
      x"FF812A01",
      x"FF7D2501",
      x"FF832B02",
      x"FF842D01",
      x"FF802703",
      x"FF802803",
      x"FF7D2500",
      x"FF872E02",
      x"FF842B01",
      x"FF862A01",
      x"FF872B01",
      x"FF882D02",
      x"FF882C02",
      x"FF892E02",
      x"FF862B00",
      x"FF8A2F02",
      x"FF8A2F00",
      x"FF8A2F02",
      x"FF892E01",
      x"FF8A2F02",
      x"FF8A2F02",
      x"FF8A2F02",
      x"FF8B3002",
      x"FF8C3200",
      x"FF8F3502",
      x"FF8D3301",
      x"FF8F3301",
      x"FF882D00",
      x"FF812803",
      x"FF7A2402",
      x"FF7D2803",
      x"FF7D2501",
      x"FF812904",
      x"FF7F2703",
      x"FF7D2801",
      x"FF7D2801",
      x"FF822A02",
      x"FF7F2802",
      x"FF802701",
      x"FF842B01",
      x"FF7F2702",
      x"FF802801",
      x"FF852C02",
      x"FF842B02",
      x"FF7E2601",
      x"FF792301",
      x"FF772301",
      x"FF772301",
      x"FF792400",
      x"FF822A01",
      x"FF7B2701",
      x"FF7F2C01",
      x"FF802901",
      x"FF7A2501",
      x"FF7E2902",
      x"FF7D2801",
      x"FF7E2901",
      x"FF7B2602",
      x"FF7C2702",
      x"FF822A03",
      x"FF802901",
      x"FF7C2702",
      x"FF802A02",
      x"FF832C01",
      x"FF7F2602",
      x"FF7D2402",
      x"FF7D2501",
      x"FF862D02",
      x"FF832A01",
      x"FF872B02",
      x"FF852A01",
      x"FF882D02",
      x"FF882C01",
      x"FF892E02",
      x"FF862B00",
      x"FF8A2F02",
      x"FF8A2F00",
      x"FF892E01",
      x"FF882D00",
      x"FF892E01",
      x"FF892E01",
      x"FF892E01",
      x"FF8B3002",
      x"FF8C3200",
      x"FF8D3301",
      x"FF8C3200",
      x"FF8E3201",
      x"FF882D00",
      x"FF802601",
      x"FF7B2301",
      x"FF7E2602",
      x"FF7B2601",
      x"FF7F2A04",
      x"FF7F2703",
      x"FF7E2902",
      x"FF7D2802",
      x"FF812901",
      x"FF822702",
      x"FF822701",
      x"FF832B01",
      x"FF7D2702",
      x"FF802803",
      x"FF832A01",
      x"FF832A01",
      x"FF7F2701",
      x"FF792301",
      x"FF772300",
      x"FF792501",
      x"FF7A2500",
      x"FF832B01",
      x"FF7C2701",
      x"FF802C01",
      x"FF802C01",
      x"FF7E2903",
      x"FF7E2903",
      x"FF7C2701",
      x"FF7C2701",
      x"FF792501",
      x"FF7C2702",
      x"FF7F2A02",
      x"FF802902",
      x"FF7F2A02",
      x"FF802B02",
      x"FF812C01",
      x"FF7B2601",
      x"FF7A2501",
      x"FF7D2501",
      x"FF852C02",
      x"FF862A01",
      x"FF872B00",
      x"FF842B01",
      x"FF852D01",
      x"FF862F01",
      x"FF882D01",
      x"FF862B00",
      x"FF892E01",
      x"FF8A2F01",
      x"FF8A2F00",
      x"FF882D00",
      x"FF882D00",
      x"FF882D01",
      x"FF892E01",
      x"FF8D3302",
      x"FF8B3001",
      x"FF8D3300",
      x"FF8C3301",
      x"FF8E3402",
      x"FF882E01",
      x"FF802702",
      x"FF792301",
      x"FF7E2901",
      x"FF802801",
      x"FF802802",
      x"FF7B2601",
      x"FF7E2902",
      x"FF7F2701",
      x"FF7F2700",
      x"FF7E2602",
      x"FF812800",
      x"FF842B03",
      x"FF7E2600",
      x"FF7F2700",
      x"FF812801",
      x"FF812801",
      x"FF7E2702",
      x"FF772402",
      x"FF782400",
      x"FF792501",
      x"FF7A2500",
      x"FF842C01",
      x"FF7C2701",
      x"FF7E2A00",
      x"FF7E2A00",
      x"FF7F2A03",
      x"FF7D2802",
      x"FF7B2600",
      x"FF7C2701",
      x"FF792601",
      x"FF7C2903",
      x"FF7E2B02",
      x"FF7E2A01",
      x"FF812801",
      x"FF832A01",
      x"FF883102",
      x"FF822A01",
      x"FF7E2803",
      x"FF7D2501",
      x"FF842B02",
      x"FF862A01",
      x"FF852C01",
      x"FF842B01",
      x"FF852D01",
      x"FF862E01",
      x"FF882D01",
      x"FF862B00",
      x"FF8A2F02",
      x"FF8B3002",
      x"FF8A2F00",
      x"FF8A2F02",
      x"FF892E01",
      x"FF872C00",
      x"FF8A2F02",
      x"FF8D3201",
      x"FF8A3000",
      x"FF8E3400",
      x"FF8D3300",
      x"FF8E3402",
      x"FF892F01",
      x"FF802803",
      x"FF792300",
      x"FF7E2903",
      x"FF7E2601",
      x"FF812900",
      x"FF7B2601",
      x"FF7E2902",
      x"FF7E2601",
      x"FF812901",
      x"FF7D2801",
      x"FF7E2600",
      x"FF832B03",
      x"FF7E2902",
      x"FF812901",
      x"FF842B03",
      x"FF812701",
      x"FF7E2702",
      x"FF772301",
      x"FF772300",
      x"FF7A2502",
      x"FF7A2500",
      x"FF842C01",
      x"FF7C2701",
      x"FF802C01",
      x"FF802B02",
      x"FF7E2903",
      x"FF7C2701",
      x"FF7B2601",
      x"FF7C2701",
      x"FF782500",
      x"FF7B2801",
      x"FF7E2A02",
      x"FF7F2B02",
      x"FF822A02",
      x"FF852C02",
      x"FF893102",
      x"FF812800",
      x"FF7C2702",
      x"FF7D2502",
      x"FF852C02",
      x"FF842900",
      x"FF842B02",
      x"FF822901",
      x"FF852C02",
      x"FF862D00",
      x"FF872C01",
      x"FF862B00",
      x"FF8A2F02",
      x"FF8A2F01",
      x"FF8A2F01",
      x"FF892E01",
      x"FF882D00",
      x"FF892E02",
      x"FF882D01",
      x"FF8D3201",
      x"FF8A2F00",
      x"FF8F3501",
      x"FF8D3200",
      x"FF8E3201",
      x"FF892F01",
      x"FF7D2701",
      x"FF782300",
      x"FF7D2802",
      x"FF7D2501",
      x"FF812901",
      x"FF7C2702",
      x"FF7F2A03",
      x"FF802802",
      x"FF802800",
      x"FF7C2701",
      x"FF7F2701",
      x"FF832B03",
      x"FF7E2902",
      x"FF802801",
      x"FF832A02",
      x"FF812802",
      x"FF7E2601",
      x"FF782302",
      x"FF772200",
      x"FF7B2502",
      x"FF7B2501",
      x"FF852E02",
      x"FF7D2801",
      x"FF802B01",
      x"FF802B03",
      x"FF7D2802",
      x"FF7C2701",
      x"FF7B2601",
      x"FF7C2702",
      x"FF7B2702",
      x"FF7C2702",
      x"FF802A02",
      x"FF802A02",
      x"FF822B02",
      x"FF832C01",
      x"FF842E01",
      x"FF802801",
      x"FF7B2501",
      x"FF7D2502",
      x"FF832A01",
      x"FF842900",
      x"FF842C02",
      x"FF822801",
      x"FF842A02",
      x"FF872C01",
      x"FF882D01",
      x"FF862B00",
      x"FF882D01",
      x"FF8A2F01",
      x"FF892E00",
      x"FF8A2F02",
      x"FF882D00",
      x"FF892E02",
      x"FF882D01",
      x"FF8D3201",
      x"FF8C3102",
      x"FF8F3501",
      x"FF8E3201",
      x"FF8E3201",
      x"FF882F01",
      x"FF7C2601",
      x"FF792202",
      x"FF7D2802",
      x"FF7E2601",
      x"FF7C2401",
      x"FF7C2702",
      x"FF7E2902",
      x"FF812903",
      x"FF7F2700",
      x"FF7F2702",
      x"FF822901",
      x"FF822902",
      x"FF802802",
      x"FF812901",
      x"FF822901",
      x"FF812802",
      x"FF7E2601",
      x"FF782302",
      x"FF782200",
      x"FF7C2603",
      x"FF7E2601",
      x"FF872F02",
      x"FF7B2701",
      x"FF7D2902",
      x"FF812B02",
      x"FF7C2702",
      x"FF7C2803",
      x"FF7B2601",
      x"FF7D2501",
      x"FF792301",
      x"FF7C2602",
      x"FF812902",
      x"FF802900",
      x"FF842C01",
      x"FF822A02",
      x"FF852D00",
      x"FF842901",
      x"FF7E2402",
      x"FF7F2502",
      x"FF842B03",
      x"FF842B01",
      x"FF802900",
      x"FF802803",
      x"FF812801",
      x"FF842B00",
      x"FF872C00",
      x"FF872C00",
      x"FF892E01",
      x"FF8A2F02",
      x"FF8A2F03",
      x"FF892E02",
      x"FF882D01",
      x"FF882D01",
      x"FF892E01",
      x"FF8C3102",
      x"FF8B3001",
      x"FF8D3301",
      x"FF8C3201",
      x"FF8C3201",
      x"FF873002",
      x"FF7C2502",
      x"FF7A2403",
      x"FF7C2603",
      x"FF792300",
      x"FF7B2601",
      x"FF7B2601",
      x"FF7C2600",
      x"FF7E2801",
      x"FF7B2601",
      x"FF7B2601",
      x"FF802601",
      x"FF7F2802",
      x"FF7F2801",
      x"FF822901",
      x"FF822901",
      x"FF812902",
      x"FF7E2602",
      x"FF7A2401",
      x"FF7A2400",
      x"FF7E2602",
      x"FF7D2501",
      x"FF8B3002",
      x"FF7C2801",
      x"FF7C2701",
      x"FF812A02",
      x"FF7B2601",
      x"FF7A2601",
      x"FF7C2702",
      x"FF7E2602",
      x"FF792301",
      x"FF7C2602",
      x"FF802903",
      x"FF802801",
      x"FF812D01",
      x"FF802A02",
      x"FF852E01",
      x"FF832B02",
      x"FF812703",
      x"FF822803",
      x"FF852D02",
      x"FF842B01",
      x"FF802900",
      x"FF802802",
      x"FF832903",
      x"FF852C01",
      x"FF882D01",
      x"FF872C01",
      x"FF892E01",
      x"FF892E01",
      x"FF892E02",
      x"FF892E02",
      x"FF872C01",
      x"FF872C01",
      x"FF882D01",
      x"FF8B3002",
      x"FF8A2F00",
      x"FF8D3301",
      x"FF8D3301",
      x"FF8D3301",
      x"FF883002",
      x"FF7A2300",
      x"FF782201",
      x"FF782201",
      x"FF7B2503",
      x"FF7B2601",
      x"FF7C2702",
      x"FF7F2902",
      x"FF7E2801",
      x"FF7B2702",
      x"FF7D2904",
      x"FF802802",
      x"FF7C2801",
      x"FF7C2800",
      x"FF832A01",
      x"FF832A01",
      x"FF822A03",
      x"FF7C2401",
      x"FF782200",
      x"FF772101",
      x"FF7E2502",
      x"FF7F2702",
      x"FF8B3102"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
