library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity img_white_mister_60 is
   port
   (
      clk       : in std_logic;
      address   : in integer range 0 to 3599; 
      data      : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of img_white_mister_60 is

   type t_rom is array(0 to 3599) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFD7D7D8",
      x"FF585959",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF484849",
      x"FFC1C1C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF959595",
      x"FFF0F1F1",
      x"FFD8D8D8",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFCFD0D0",
      x"FFF7F7F8",
      x"FF747575",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF575858",
      x"FFD6D7D7",
      x"FF141414",
      x"FF646464",
      x"FFC8C8C8",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFAFAFB0",
      x"FF707070",
      x"FF131313",
      x"FFC7C8C8",
      x"FF383939",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC8C9C9",
      x"FF707171",
      x"FF000000",
      x"FF040404",
      x"FFAEAEAF",
      x"FF929292",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF6C6C6D",
      x"FFAFAFB0",
      x"FF060707",
      x"FF000000",
      x"FF747474",
      x"FF989999",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF5C5D5D",
      x"FFC2C2C2",
      x"FF19191A",
      x"FF92476E",
      x"FF673552",
      x"FF272728",
      x"FFD0D0D1",
      x"FF545455",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFD6D6D6",
      x"FF2D2D2D",
      x"FF64334F",
      x"FF984973",
      x"FF1C1B1B",
      x"FFC4C4C4",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9BABA",
      x"FF747576",
      x"FF090407",
      x"FFB65889",
      x"FFA5507E",
      x"FF070305",
      x"FF616162",
      x"FFCECECE",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB0B0B1",
      x"FF6A6A6A",
      x"FF060305",
      x"FFA04F7B",
      x"FFB8598B",
      x"FF0B0507",
      x"FF7B7B7C",
      x"FF949495",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF626262",
      x"FFF5F5F6",
      x"FF181818",
      x"FF0B0B0B",
      x"FF171717",
      x"FF181918",
      x"FF101010",
      x"FF0C0C0C",
      x"FFD3D4D5",
      x"FFACADAD",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF848384",
      x"FFDCDDDD",
      x"FF0D0D0D",
      x"FF101010",
      x"FF181818",
      x"FF171717",
      x"FF0B0B0B",
      x"FF131313",
      x"FFDEDEDE",
      x"FF363636",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC8C9CA",
      x"FFF1F2F3",
      x"FFAFB0B1",
      x"FFAAABAB",
      x"FFC1C1C1",
      x"FFC2C3C2",
      x"FFB3B4B5",
      x"FFABACAD",
      x"FFE7E8E9",
      x"FFF4F5F6",
      x"FF868788",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF737475",
      x"FF787979",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFACADAD",
      x"FFB3B4B5",
      x"FFC2C2C2",
      x"FFC1C1C1",
      x"FFABACAC",
      x"FFAEAFAF",
      x"FFF2F3F3",
      x"FF838383",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFAFAFAF",
      x"FFF3F3F3",
      x"FFEEEFF0",
      x"FFE5E6E7",
      x"FFEDEEEF",
      x"FFEDEEEF",
      x"FFE9EAEB",
      x"FFE8E9EA",
      x"FFECEDEE",
      x"FFEDEEEF",
      x"FFE6E7E8",
      x"FFE5E6E7",
      x"FFF6F6F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFEDEEEF",
      x"FFECEDEE",
      x"FFE8EAEB",
      x"FFE9EAEB",
      x"FFEDEEEF",
      x"FFEDEEEF",
      x"FFE7E8E9",
      x"FFEDEEEE",
      x"FFB8B9B9",
      x"FF5E5E5E",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA6A7A7",
      x"FFF2F3F4",
      x"FFE9EAEB",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFEEEFF0",
      x"FFEDEDEE",
      x"FF747575",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF737374",
      x"FFF5F6F6",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFEBEBEC",
      x"FF525253",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB1B1B2",
      x"FFEEEFF0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF0F0F1",
      x"FF9D9D9D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBDBDBE",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFC2C3C3",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBABBBB",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFC2C2C3",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9B9BA",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFC2C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9B9BA",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFC2C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9B9BA",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEBECED",
      x"FFE8E9E9",
      x"FFE8E9E9",
      x"FFEBECED",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEBECED",
      x"FFE7E8E8",
      x"FFE9E9EA",
      x"FFEAECEC",
      x"FFE6E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFC2C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9B9BA",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEBECED",
      x"FFE1E1E2",
      x"FF444545",
      x"FF424343",
      x"FFDFE0E1",
      x"FFEBECED",
      x"FFEBECED",
      x"FFDBDBDC",
      x"FF3E3F3F",
      x"FF494949",
      x"FFE5E5E6",
      x"FFEAEBEC",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFC2C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9B9BA",
      x"FFF4F4F5",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFEFF0F2",
      x"FFF4F5F6",
      x"FF959596",
      x"FF000000",
      x"FF000000",
      x"FF848585",
      x"FFF2F3F4",
      x"FFF5F5F6",
      x"FF838383",
      x"FF000000",
      x"FF000000",
      x"FF9E9F9F",
      x"FFF5F6F6",
      x"FFF0F1F2",
      x"FFF0F1F2",
      x"FFF0F1F2",
      x"FFF0F1F2",
      x"FFF0F1F1",
      x"FFEFF0F1",
      x"FFF0F1F2",
      x"FFF0F1F2",
      x"FFEFF0F1",
      x"FFEFF0F2",
      x"FFF0F1F2",
      x"FFEFF0F1",
      x"FFEFF0F1",
      x"FFEFF0F2",
      x"FFF4F4F5",
      x"FFC2C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB9B9BA",
      x"FFB6B6B7",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5A5A5A",
      x"FF5D5D5E",
      x"FF3E3F3F",
      x"FF000000",
      x"FF000000",
      x"FF212121",
      x"FF686868",
      x"FF717171",
      x"FF282929",
      x"FF000000",
      x"FF000000",
      x"FF474848",
      x"FF686868",
      x"FF636364",
      x"FF636364",
      x"FF616263",
      x"FF616263",
      x"FF606161",
      x"FF606061",
      x"FF5E5F60",
      x"FF5E5F5F",
      x"FF5D5E5E",
      x"FF5D5D5D",
      x"FF5C5C5C",
      x"FF5B5C5C",
      x"FF5A5B5B",
      x"FF5A5A5A",
      x"FFBBBBBC",
      x"FFC1C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC3C4C4",
      x"FF5B5B5B",
      x"FF010101",
      x"FF050505",
      x"FF060606",
      x"FF060606",
      x"FF060606",
      x"FF060606",
      x"FF040404",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF040404",
      x"FF060606",
      x"FF060606",
      x"FF060606",
      x"FF050505",
      x"FF010101",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF010101",
      x"FF020202",
      x"FF020202",
      x"FF030303",
      x"FF020202",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF030303",
      x"FF050505",
      x"FF050505",
      x"FF050505",
      x"FF050505",
      x"FF040404",
      x"FF000000",
      x"FF606061",
      x"FFC9C9CA",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC5C6C6",
      x"FF4D4E4E",
      x"FF0F0F0F",
      x"FF808080",
      x"FFAAAAAA",
      x"FFAAAAAA",
      x"FFAAAAAA",
      x"FFAAAAAA",
      x"FF787878",
      x"FF060606",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF7E7E7E",
      x"FFAAAAAA",
      x"FFAAAAAA",
      x"FFAAAAAA",
      x"FF9A9A9A",
      x"FF292929",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF262626",
      x"FF8E8E8E",
      x"FF9E9E9E",
      x"FF9E9E9E",
      x"FF9F9F9F",
      x"FF717171",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF090909",
      x"FF767676",
      x"FFA6A6A6",
      x"FFA7A7A7",
      x"FFA8A8A8",
      x"FFA9A9A9",
      x"FF7F7F7F",
      x"FF0C0C0C",
      x"FF505050",
      x"FFCCCCCD",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC7C8C8",
      x"FF535454",
      x"FF101010",
      x"FFB9B9B9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCDCDCD",
      x"FF232323",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF111111",
      x"FFEBEBEB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE7E7E7",
      x"FF3D3D3D",
      x"FF0F0F0F",
      x"FF606063",
      x"FF5B5B5E",
      x"FF0C0C0D",
      x"FF434343",
      x"FFEDEDED",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFE7E7E7",
      x"FF0E0E0E",
      x"FF000000",
      x"FF000000",
      x"FF000000",
      x"FF272727",
      x"FFD1D1D1",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFB4B4B4",
      x"FF0B0B0B",
      x"FF565656",
      x"FFCCCCCC",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBCBCBD",
      x"FF6B6C6B",
      x"FF020202",
      x"FF939393",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF8F8F8",
      x"FF989898",
      x"FF0B0B0B",
      x"FF000000",
      x"FF141414",
      x"FF969696",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCCCCCC",
      x"FF222222",
      x"FF1F1F20",
      x"FF949599",
      x"FF939497",
      x"FF1D1D1E",
      x"FF272727",
      x"FFD1D1D1",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF8F8F8F",
      x"FF121212",
      x"FF000000",
      x"FF0D0D0D",
      x"FF9E9E9E",
      x"FFF9F9F9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF888888",
      x"FF010101",
      x"FF717272",
      x"FFC3C3C4",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF595A5A",
      x"FFDFE0E0",
      x"FFAFAFB0",
      x"FF000000",
      x"FF2B2B2B",
      x"FFFBFBFB",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFECECEC",
      x"FFCBCBCB",
      x"FFEEEEEE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FF878787",
      x"FF010101",
      x"FF121213",
      x"FF313132",
      x"FF2F2F30",
      x"FF0F0F0F",
      x"FF030303",
      x"FF8E8E8E",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFECECEC",
      x"FFCCCCCC",
      x"FFEEEEEE",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF8F8F8",
      x"FF252525",
      x"FF000000",
      x"FFB6B7B8",
      x"FFEFF0F0",
      x"FF8A8A8A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC7C7C7",
      x"FFEEEFEF",
      x"FFEDEEEF",
      x"FFEDEDEE",
      x"FF1D1D1D",
      x"FF000000",
      x"FFA9A9A9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFCDCDCD",
      x"FF191919",
      x"FF000000",
      x"FF000000",
      x"FF010101",
      x"FF010101",
      x"FF000000",
      x"FF000000",
      x"FF1B1B1B",
      x"FF9A9A9A",
      x"FFF2F2F2",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFA0A0A0",
      x"FF010101",
      x"FF232324",
      x"FFEEEFF0",
      x"FFEBECED",
      x"FFEFEFF0",
      x"FFD0D0D0",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF393939",
      x"FFDADADA",
      x"FFEEEFF0",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFF1F2F3",
      x"FFA2A2A3",
      x"FF0E0E0E",
      x"FF1C1C1C",
      x"FFAAAAAA",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF5F5F5",
      x"FF757575",
      x"FF0F0F0F",
      x"FF161616",
      x"FF020102",
      x"FF974269",
      x"FFE369A7",
      x"FFE369A7",
      x"FFA54974",
      x"FF0B0408",
      x"FF1B1B1C",
      x"FF161616",
      x"FF343434",
      x"FFD8D8D8",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFA5A5A5",
      x"FF191919",
      x"FF0F0F0F",
      x"FFA8A8A8",
      x"FFEFF0F1",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFEEEFF0",
      x"FFD7D8D8",
      x"FF343535",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFABACAC",
      x"FFF2F2F3",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFE9E9EA",
      x"FF6D6D6E",
      x"FF000000",
      x"FF1D1D1D",
      x"FFAAAAAA",
      x"FFF8F8F8",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF8F8F8",
      x"FF818181",
      x"FF0A0A0A",
      x"FF5D5E5E",
      x"FF919293",
      x"FF0B0B0B",
      x"FF210E17",
      x"FF853F64",
      x"FF874066",
      x"FF230F19",
      x"FF050404",
      x"FF7E7E80",
      x"FFA0A0A2",
      x"FF1D1D1E",
      x"FF424242",
      x"FFD9D9D9",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFFFFFFF",
      x"FFF6F6F6",
      x"FFA5A5A5",
      x"FF1B1B1B",
      x"FF000000",
      x"FF747474",
      x"FFEAEAEB",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFF2F3F3",
      x"FFA9AAAA",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFF9F9F9",
      x"FFE9EAEB",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFF8F8F9",
      x"FF6F6F6F",
      x"FF0F0F0F",
      x"FF010101",
      x"FF363636",
      x"FF9B9B9B",
      x"FFC5C5C5",
      x"FFD7D7D7",
      x"FFD9D9D9",
      x"FFCCCCCC",
      x"FFB3B3B3",
      x"FF535353",
      x"FF070707",
      x"FF666667",
      x"FFC9C9CC",
      x"FFC1C2C4",
      x"FFBFC0C1",
      x"FF4B4B4B",
      x"FF080909",
      x"FF070807",
      x"FF454546",
      x"FFB9BABC",
      x"FFC0C1C3",
      x"FFC6C7C9",
      x"FFA1A2A4",
      x"FF111111",
      x"FF3E3E3E",
      x"FFB5B5B5",
      x"FFCDCDCD",
      x"FFD9D9D9",
      x"FFD7D7D7",
      x"FFC4C4C4",
      x"FF999999",
      x"FF323232",
      x"FF000000",
      x"FF101010",
      x"FF747575",
      x"FFF6F6F7",
      x"FFE8E9EA",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE8E9EA",
      x"FFF8F9F9",
      x"FF363636",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF606061",
      x"FFF7F7F7",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFEBECEC",
      x"FFA0A0A0",
      x"FF202020",
      x"FF000000",
      x"FF050505",
      x"FF1B1B1B",
      x"FF2D2D2D",
      x"FF2F2F2F",
      x"FF222222",
      x"FF0D0D0D",
      x"FF000000",
      x"FF010101",
      x"FF2F2F2F",
      x"FFA4A5A7",
      x"FFC0C1C3",
      x"FFC8C9CB",
      x"FFB5B6B8",
      x"FF929495",
      x"FF909193",
      x"FFB1B2B4",
      x"FFC9CACC",
      x"FFBDBEC0",
      x"FFC0C1C3",
      x"FF4E4F50",
      x"FF080808",
      x"FF000000",
      x"FF0E0E0E",
      x"FF232323",
      x"FF2F2F2F",
      x"FF2D2D2D",
      x"FF1A1A1A",
      x"FF050505",
      x"FF000000",
      x"FF232323",
      x"FFA3A3A3",
      x"FFEBEBEC",
      x"FFE8EAEB",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF6F7F7",
      x"FF747475",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF79797A",
      x"FFF7F7F8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFF1F2F2",
      x"FFECECED",
      x"FFABABAB",
      x"FF575656",
      x"FF373737",
      x"FF292929",
      x"FF272727",
      x"FF303030",
      x"FF0A0A0A",
      x"FF000000",
      x"FF616162",
      x"FFC5C6C6",
      x"FF828384",
      x"FFC7C8CA",
      x"FFC5C6C8",
      x"FFCBCCCE",
      x"FF7E7F80",
      x"FF7B7B7C",
      x"FFCECFD1",
      x"FFC1C2C4",
      x"FFC5C6C8",
      x"FF969798",
      x"FFA7A8AA",
      x"FF939395",
      x"FF0B0B0B",
      x"FF020303",
      x"FF252525",
      x"FF292929",
      x"FF292929",
      x"FF373838",
      x"FF585858",
      x"FFADAEAF",
      x"FFECEDED",
      x"FFF1F2F2",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF5F6F7",
      x"FF919192",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF777777",
      x"FFF7F7F8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFEAEBEC",
      x"FFEFF0F0",
      x"FFEEEEEF",
      x"FFE1E1E1",
      x"FFD3D3D3",
      x"FFD1D1D1",
      x"FFA2A2A2",
      x"FF494949",
      x"FF373838",
      x"FF2B2B2C",
      x"FF3A3B3B",
      x"FF868789",
      x"FFD8D9DB",
      x"FFB7B8B9",
      x"FF575758",
      x"FF0E0E0E",
      x"FF101010",
      x"FF6E6F70",
      x"FFC3C4C6",
      x"FFD5D6D9",
      x"FFABACAE",
      x"FF333333",
      x"FF2B2B2B",
      x"FF282828",
      x"FF616162",
      x"FF606060",
      x"FFD3D3D3",
      x"FFD3D3D3",
      x"FFE1E2E2",
      x"FFEEEFEF",
      x"FFEFF0F0",
      x"FFEAEBEC",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF6F7F7",
      x"FF8E8E8F",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF4C4C4D",
      x"FFF7F7F8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEBECED",
      x"FFEBECED",
      x"FF252525",
      x"FFC1C1C1",
      x"FFA6A6A6",
      x"FF111111",
      x"FF0F0F0F",
      x"FF343535",
      x"FF1F2020",
      x"FF090909",
      x"FF1F1F20",
      x"FF1E1E1F",
      x"FF1D1D1E",
      x"FF171718",
      x"FF0A0A0B",
      x"FF272728",
      x"FF2C2C2D",
      x"FF0F0F0F",
      x"FF171717",
      x"FF747474",
      x"FFE5E5E5",
      x"FF3D3D3E",
      x"FFB8B9B9",
      x"FFEEEFEF",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF6F7F7",
      x"FF666666",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFE3E4E4",
      x"FFEBECED",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFA0A1A1",
      x"FF4E4F4F",
      x"FFF6F6F6",
      x"FF414141",
      x"FF828282",
      x"FF818282",
      x"FF444445",
      x"FF000000",
      x"FF0E0E0E",
      x"FF636467",
      x"FF77777A",
      x"FF77787C",
      x"FF5D5D60",
      x"FF0A0A0A",
      x"FF000000",
      x"FF383838",
      x"FF868787",
      x"FFABACAC",
      x"FF393939",
      x"FFE7E8E8",
      x"FF8E8E8E",
      x"FF5A5B5B",
      x"FFF0F1F1",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEBECED",
      x"FFF3F3F3",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF5A5A5A",
      x"FFE9EAEB",
      x"FFE9EAEB",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF2F2F3",
      x"FF5B5B5C",
      x"FF8A8A8A",
      x"FFC7C7C8",
      x"FF404041",
      x"FFE7E8E9",
      x"FFF6F7F8",
      x"FFF9F9FA",
      x"FF8D8E8E",
      x"FF3B3B3B",
      x"FF141414",
      x"FF040404",
      x"FF030303",
      x"FF111111",
      x"FF333333",
      x"FF7D7D7D",
      x"FFF4F5F5",
      x"FFF5F6F7",
      x"FFF4F4F5",
      x"FF6D6D6D",
      x"FF727272",
      x"FFE1E2E3",
      x"FF363636",
      x"FFDFDFE0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE8E9EA",
      x"FFEBEBEC",
      x"FF727273",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF717171",
      x"FFFBFBFB",
      x"FFEDEEEF",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFF0F1F1",
      x"FF818282",
      x"FFAFAFB0",
      x"FF7E7F7F",
      x"FF656666",
      x"FFF1F2F2",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFEFEFF1",
      x"FFE1E1E1",
      x"FFBABABA",
      x"FF9A9A9B",
      x"FF979898",
      x"FFB6B6B6",
      x"FFDDDDDD",
      x"FFEFF0F0",
      x"FFEAEBEC",
      x"FFE7E8E9",
      x"FFEEEFF0",
      x"FFB4B5B5",
      x"FF4B4C4C",
      x"FFECECED",
      x"FF646566",
      x"FFDEDFE0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFEBECED",
      x"FFF8F9F9",
      x"FF8B8B8B",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF404141",
      x"FFACACAC",
      x"FFE9EAEB",
      x"FFE8E9EA",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFF1F2F3",
      x"FFFBFBFB",
      x"FF5C5C5C",
      x"FF858585",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEAEBED",
      x"FFF1F2F3",
      x"FFF2F3F4",
      x"FFECEDEE",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFD7D8D9",
      x"FF383839",
      x"FFE2E2E2",
      x"FFF4F5F6",
      x"FFE8E9EA",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEAEBEB",
      x"FFBBBBBB",
      x"FF5A5A5B",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBEBEC0",
      x"FFEEEFEF",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEDEEEF",
      x"FFA3A4A5",
      x"FFB4B5B5",
      x"FFEBECED",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEBEBEC",
      x"FFDFDFE0",
      x"FF909192",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEEEEEF",
      x"FFC1C2C2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBBBCBD",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFF1F1F2",
      x"FFF0F1F2",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFE8E9EA",
      x"FFF3F3F4",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFBABBBB",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBBBCBD",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFBBBCBC",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBBBCBD",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFBBBCBC",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBBBCBD",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFBBBCBC",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBBBCBD",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFBABBBB",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFB5B6B7",
      x"FFEFF0F0",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEFF0F0",
      x"FFB8B9B9",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF414142",
      x"FF7A7A7A",
      x"FFDADADB",
      x"FFEAEBEC",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEDEEEF",
      x"FFF1F1F2",
      x"FFF1F2F3",
      x"FFF1F2F3",
      x"FFF1F1F2",
      x"FFEEEFEF",
      x"FFE8E9EA",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE8E9EA",
      x"FFE6E7E8",
      x"FFA5A5A5",
      x"FF4A4A4A",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF474748",
      x"FFE3E3E4",
      x"FFF2F3F4",
      x"FFE9EAEB",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E8E9",
      x"FFE8EAEB",
      x"FFF5F6F6",
      x"FFD4D4D4",
      x"FF929293",
      x"FF777777",
      x"FF777777",
      x"FF919191",
      x"FFD1D2D3",
      x"FFF4F5F6",
      x"FFE9EAEB",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFF0F1F1",
      x"FFE4E4E4",
      x"FF4C4D4D",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFC2C2C2",
      x"FFEAEBEC",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFEFF1F1",
      x"FFD9D9D9",
      x"FF505050",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF4C4C4D",
      x"FFD6D6D7",
      x"FFF0F1F2",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E9EA",
      x"FFD1D2D2",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFD0D1D1",
      x"FFE6E7E8",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFEAEBEC",
      x"FFD6D6D6",
      x"FF414141",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF3D3D3D",
      x"FFD4D4D4",
      x"FFEBECED",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE6E7E8",
      x"FFE8E9E9",
      x"FF3F4040",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFBABABB",
      x"FFECEDED",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE9EAEB",
      x"FFEFF0F0",
      x"FF353535",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFEEEEEE",
      x"FFEAEBEC",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFE7E8E9",
      x"FFDBDBDB",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF565857",
      x"FFFCFCFC",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF9F9F9",
      x"FFACACAC",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FFA5A5A5",
      x"FFFAFAFA",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF7F7F8",
      x"FFF8F8F8",
      x"FF8B8B8C",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF4B4B4B",
      x"FF848484",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF848586",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"FF848585",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF808181",
      x"FF828384",
      x"FF5A5B5B",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(address);
      end if;
   end process;

end architecture;
